library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.common.all;
use work.rendering_common.all;

entity renderer_triangle is
	port(
		clk           : in  std_logic;
		rst           : in  std_logic;
		tile_rect_in  : in  rect_t;
		triangle_in   : in  triangle2d_t;
		put_pixel_out : out std_logic;
		posx_out      : out unsigned(15 downto 0);
		posy_out      : out unsigned(15 downto 0);
		start_in      : in  std_logic;
		ready_out     : out std_logic;
		area_in       : in  int32_t;
		depths_in     : in  point3d_t;
		colors_in     : in  triangle_colors_t;
		color_out     : out color_t;
		depth_buf_in : out unsigned(15 downto 0);
		depth_buf_out : in unsigned(15 downto 0);
		depth_wren : out std_logic
	);
end entity renderer_triangle;

architecture RTL of renderer_triangle is

	-- BOUNDING BOX CALCULATION

	signal render_rect_latch, render_rect_latch_next : srect_t;

	

	signal depth_out_latch : unsigned(15 downto 0);

	-- TRIANGLE RENDERING

	signal cntx, cntx_next : int16_t := (others => '0');
	signal cnty, cnty_next : int16_t := (others => '0');

	signal put_pixel_out_next : std_logic := '0';
	signal ready_out_next     : std_logic := '0';

	signal triangle_latch, triangle_latch_next : triangle2d_t := (point2d(0, 0), point2d(0, 0), point2d(0, 0));

	function cross_product(x, y : int16_t; p2, p3 : point2d_t) return int32_t is
	begin
		return ((x - p3.x) * (p2.y - p3.y) - (p2.x - p3.x) * (y - p3.y));
	end function;
	
	function interpolate_color_component(
		c0, c1, c2 : std_logic_vector(7 downto 0);
		e0, e1, e2 : int32_t;
		area : int32_t
	) return int32_t is
	begin
		return resize(
				e0 * signed('0' & c0) + 
				e1 * signed('0' & c1) + 
				e2 * signed('0' & c2), 32
		) / area;
	end function;

	-- CONTROL

	type state_type is (
		st_start, st_idle, st_render, st_finished, st_start_render, st_wait_0
	);
	signal state, state_next : state_type := st_start;

begin
	posx_out <= uint16_with_cut(cntx);
	posy_out <= uint16_with_cut(cnty);

	process(clk, rst) is
	begin
		if rst = '1' then
			state <= st_start;
		elsif rising_edge(clk) then
			put_pixel_out     <= put_pixel_out_next;
			cntx              <= cntx_next;
			cnty              <= cnty_next;
			ready_out         <= ready_out_next;
			render_rect_latch <= render_rect_latch_next;
			state             <= state_next;
			triangle_latch    <= triangle_latch_next;
		end if;
	end process;

	process(state, cntx, cnty, render_rect_latch.x0, render_rect_latch.x1, render_rect_latch.y0, render_rect_latch.y1, put_pixel_out, ready_out, start_in, render_rect_latch, tile_rect_in, triangle_in, triangle_latch, area_in, depths_in.x, depths_in.y, depths_in.z, colors_in(0).b, colors_in(0).g, colors_in(0).r, colors_in(1).r, colors_in(2).r, colors_in(1).b, colors_in(1).g, colors_in(2).b, colors_in(2).g, depth_buf_out, depth_out_latch) is
		variable e0, e1, e2 : int32_t;
		variable depth      : signed(47 downto 0);
		variable r, g, b : int32_t;
	begin
		state_next             <= state;
		put_pixel_out_next     <= put_pixel_out;
		cntx_next              <= cntx;
		cnty_next              <= cnty;
		ready_out_next         <= ready_out;
		render_rect_latch_next <= render_rect_latch;
		triangle_latch_next    <= triangle_latch;

		case state is
		when st_start =>
				depth_wren <= '0';
				put_pixel_out_next  <= '0';
				cntx_next           <= (others => '0');
				cnty_next           <= (others => '0');
				ready_out_next      <= '0';
				triangle_latch_next <= (point2d(0, 0), point2d(0, 0), point2d(0, 0));
				state_next          <= st_idle;

			when st_idle =>
				depth_wren <= '0';
				put_pixel_out_next <= '0';
				ready_out_next     <= '0';
				if start_in = '1' then
					triangle_latch_next    <= triangle_in;
					render_rect_latch_next <= get_current_rendering_bounding_box(triangle_in, tile_rect_in);
					state_next             <= st_start_render;
				else
					state_next <= st_idle;
				end if;

			when st_start_render =>
				put_pixel_out_next <= '0';
				depth_wren <= '0';
				cntx_next          <= render_rect_latch.x0;
				cnty_next          <= render_rect_latch.y0;

				state_next <= st_render;

			when st_render =>
				put_pixel_out_next <= '0';
				depth_wren <= '0';

				if cnty <= render_rect_latch.y1 then
					if cntx < render_rect_latch.x1 then
						e0 := cross_product(cntx, cnty, triangle_latch(0), triangle_latch(1));
						e1 := cross_product(cntx, cnty, triangle_latch(1), triangle_latch(2));
						e2 := cross_product(cntx, cnty, triangle_latch(2), triangle_latch(0));


						if e0 <= 0 and e1 <= 0 and e2 <= 0 then

							r := interpolate_color_component(colors_in(2).r, colors_in(0).r, colors_in(1).r, e0, e1, e2, area_in);
							g := interpolate_color_component(colors_in(2).g, colors_in(0).g, colors_in(1).g, e0, e1, e2, area_in);
							b := interpolate_color_component(colors_in(2).b, colors_in(0).b, colors_in(1).b, e0, e1, e2, area_in);
----							

							depth_out_latch <= depth_buf_out;
							depth := 256 - (e0 * depths_in.z + e1 * depths_in.x + e2 * depths_in.y) / area_in;

							state_next <= st_wait_0;
						else
							cntx_next <= cntx + 1;
						end if;

						
					else
						cntx_next <= render_rect_latch.x0;
						cnty_next <= cnty + 1;
					end if;
				else
					ready_out_next     <= '1';
					put_pixel_out_next <= '0';
					state_next         <= st_idle;
				end if;
				
			when st_wait_0 =>
				depth_wren <= '0';
				if unsigned(std_logic_vector(depth+127))(15 downto 0) > depth_out_latch then
					depth_wren <= '1';
					depth_buf_in <= unsigned(std_logic_vector(depth+127))(15 downto 0);
					--color_out <= (
					--	r => std_logic_vector(depth)(7 downto 0),
					--	g => std_logic_vector(depth)(7 downto 0),
					--	b => std_logic_vector(depth)(7 downto 0)
					--);
					color_out <= (
						r => std_logic_vector(r)(7 downto 0),
						g => std_logic_vector(g)(7 downto 0),
						b => std_logic_vector(b)(7 downto 0)
					);
--							color_out <= (
--								r => X"00",
--								g => X"5F",
--								b => X"FF"
--							);

					put_pixel_out_next <= '1';
				else
					put_pixel_out_next <= '0';
				end if;
				cntx_next <= cntx + 1;
				state_next <= st_render;
				
			when st_finished =>
				depth_wren <= '0';
				ready_out_next     <= '1';
				put_pixel_out_next <= '0';
				cntx_next          <= (others => '0');
				cnty_next          <= (others => '0');

				state_next <= st_start;
		end case;
	end process;

end architecture RTL;