use work.common.all;

package renderer_mesh is
	constant vertices : vertex_arr_3d_t(0 to 90) := (
		point3d(439, 134, 80), point3d(401, 194, 80), point3d(401, 194, 71), point3d(439, 134, 71), point3d(407, 198, 80), point3d(448, 134, 80), point3d(307, 218, 80), point3d(307, 218, 71), point3d(307, 224, 80), point3d(211, 194, 80), point3d(213, 194, 71), 
		point3d(207, 198, 80), point3d(176, 134, 80), point3d(176, 134, 71), point3d(166, 134, 80), point3d(430, 213, 151), point3d(481, 134, 151), point3d(441, 219, 217), point3d(495, 134, 217), point3d(307, 245, 151), point3d(307, 255, 217), 
		point3d(184, 213, 151), point3d(174, 219, 217), point3d(134, 134, 151), point3d(119, 134, 217), point3d(424, 209, 264), point3d(472, 134, 264), point3d(407, 198, 286), point3d(448, 134, 286), point3d(307, 239, 264), point3d(307, 224, 286), 
		point3d(191, 209, 264), point3d(207, 198, 286), point3d(143, 134, 264), point3d(166, 134, 286), point3d(393, 189, 295), point3d(428, 134, 295), point3d(307, 134, 300), point3d(307, 211, 295), point3d(222, 189, 295), point3d(187, 134, 295), 
		point3d(157, 134, 114), point3d(162, 147, 104), point3d(71, 147, 108), point3d(81, 134, 117), point3d(40, 147, 135), point3d(54, 134, 135), point3d(166, 134, 94), point3d(61, 134, 99), point3d(25, 134, 135), point3d(60, 147, 185), 
		point3d(69, 134, 176), point3d(124, 147, 231), point3d(51, 134, 194), point3d(129, 134, 245), point3d(467, 134, 169), point3d(467, 164, 207), point3d(546, 154, 151), point3d(532, 134, 135), point3d(589, 145, 80), point3d(561, 134, 80), 
		point3d(467, 134, 245), point3d(560, 134, 168), point3d(617, 134, 80), point3d(601, 143, 74), point3d(573, 134, 75), point3d(589, 140, 80), point3d(570, 134, 80), point3d(630, 134, 73), point3d(608, 134, 80), point3d(307, 134, 11), 
		point3d(329, 148, 27), point3d(338, 134, 27), point3d(321, 142, 53), point3d(326, 134, 53), point3d(307, 153, 27), point3d(307, 146, 53), point3d(286, 148, 27), point3d(294, 142, 53), point3d(277, 134, 27), point3d(289, 134, 53), 
		point3d(362, 169, 66), point3d(385, 134, 66), point3d(394, 189, 80), point3d(430, 134, 80), point3d(307, 183, 66), point3d(307, 212, 80), point3d(252, 169, 66), point3d(221, 189, 80), point3d(230, 134, 66), point3d(185, 134, 80)
		
	);

	constant indices : indices_arr_t(0 to 129) := (
		idx(0, 1, 2), idx(2, 3, 0), 
		idx(3, 2, 4), idx(4, 5, 3), idx(1, 6, 7), idx(7, 2, 1), idx(2, 7, 8), idx(8, 4, 2), idx(6, 9, 10), idx(10, 7, 6), idx(7, 10, 11), idx(11, 8, 7), 
		idx(9, 12, 13), idx(13, 10, 9), idx(10, 13, 14), idx(14, 11, 10), idx(5, 4, 15), idx(15, 16, 5), idx(16, 15, 17), idx(17, 18, 16), idx(4, 8, 19), idx(19, 15, 4), 
		idx(15, 19, 20), idx(20, 17, 15), idx(8, 11, 21), idx(21, 19, 8), idx(19, 21, 22), idx(22, 20, 19), idx(11, 14, 23), idx(23, 21, 11), idx(21, 23, 24), idx(24, 22, 21), 
		idx(18, 17, 25), idx(25, 26, 18), idx(26, 25, 27), idx(27, 28, 26), idx(17, 20, 29), idx(29, 25, 17), idx(25, 29, 30), idx(30, 27, 25), idx(20, 22, 31), idx(31, 29, 20), 
		idx(29, 31, 32), idx(32, 30, 29), idx(22, 24, 33), idx(33, 31, 22), idx(31, 33, 34), idx(34, 32, 31), idx(28, 27, 35), idx(35, 36, 28), idx(36, 35, 37), idx(37, 37, 36), 
		idx(27, 30, 38), idx(38, 35, 27), idx(35, 38, 37), idx(37, 37, 35), idx(30, 32, 39), idx(39, 38, 30), idx(38, 39, 37), idx(37, 37, 38), idx(32, 34, 40), idx(40, 39, 32), 
		idx(39, 40, 37), idx(37, 37, 39), idx(37, 37, 40), idx(41, 42, 43), idx(43, 44, 41), idx(44, 43, 45), idx(45, 46, 44), idx(42, 47, 48), idx(48, 43, 42), idx(43, 48, 49), 
		idx(49, 45, 43), idx(46, 45, 50), idx(50, 51, 46), idx(51, 50, 52), idx(52, 24, 51), idx(45, 49, 53), idx(53, 50, 45), idx(50, 53, 54), idx(54, 52, 50), idx(55, 56, 57), 
		idx(57, 58, 55), idx(58, 57, 59), idx(59, 60, 58), idx(56, 61, 62), idx(62, 57, 56), idx(57, 62, 63), idx(63, 59, 57), idx(60, 59, 64), idx(64, 65, 60), idx(65, 64, 66), 
		idx(66, 67, 65), idx(59, 63, 68), idx(68, 64, 59), idx(64, 68, 69), idx(69, 66, 64), idx(70, 70, 71), idx(71, 72, 70), idx(72, 71, 73), idx(73, 74, 72), idx(70, 70, 75), 
		idx(75, 71, 70), idx(71, 75, 76), idx(76, 73, 71), idx(70, 70, 77), idx(77, 75, 70), idx(75, 77, 78), idx(78, 76, 75), idx(70, 70, 79), idx(79, 77, 70), idx(77, 79, 80), 
		idx(80, 78, 77), idx(70, 70, 72), idx(74, 73, 81), idx(81, 82, 74), idx(82, 81, 83), idx(83, 84, 82), idx(73, 76, 85), idx(85, 81, 73), idx(81, 85, 86), idx(86, 83, 81), 
		idx(76, 78, 87), idx(87, 85, 76), idx(85, 87, 88), idx(88, 86, 85), idx(78, 80, 89), idx(89, 87, 78), idx(87, 89, 90), idx(90, 88, 87)
	);

end package renderer_mesh;
