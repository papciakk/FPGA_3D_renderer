use work.definitions.all;

package mesh is
	constant vertices : vertex_attr_arr_t(0 to 25) := (
		va(18726, -20751, -40, 14138, -29560, 0), va(12391, -20751, 15468, 9964, -29583, 9964), va(10162, -22253, 13239, 6607, -31406, 6607), 
		va(15586, -22253, -40, 9339, -31408, 0), va(-3117, -22936, -40, 0, -32767, 0), va(-3117, -20751, 21803, 0, -29560, 14138), 
		va(-3117, -22253, 18663, 0, -31408, 9339), va(-18626, -20751, 15468, -9964, -29583, 9964), va(-16397, -22253, 13239, -6607, -31406, 6607), 
		va(-24961, -20751, -40, -14138, -29560, 0), va(-21821, -22253, -40, -9339, -31408, 0), va(-18626, -20751, -15549, -9964, -29583, -9964), 
		va(-16397, -22253, -13320, -6607, -31406, -6607), va(-3117, -20751, -21884, 0, -29560, -14138), va(-3117, -22253, -18744, 0, -31408, -9339), 
		va(12391, -20751, -15549, 9964, -29583, -9964), va(10162, -22253, -13320, 6607, -31406, -6607), va(-3117, 22936, -40, 0, 32767, 0), 
		va(247, 20478, 3323, 10632, 29113, 10632), va(1615, 20478, -40, 15100, 29081, 0), va(-3117, 20478, 4692, 0, 29081, 15100), 
		va(-6481, 20478, 3323, -10632, 29113, 10632), va(-7850, 20478, -40, -15100, 29081, 0), va(-6481, 20478, -3405, -10632, 29113, -10632), 
		va(-3117, 20478, -4773, 0, 29081, -15100), va(247, 20478, -3405, 10632, 29113, -10632)
	);

	constant indices : indices_arr_t(0 to 47) := (
		idx(0, 1, 2), idx(2, 3, 0), idx(3, 2, 4), idx(4, 4, 3), idx(1, 5, 6), 
		idx(6, 2, 1), idx(2, 6, 4), idx(4, 4, 2), idx(5, 7, 8), idx(8, 6, 5), 
		idx(6, 8, 4), idx(4, 4, 6), idx(7, 9, 10), idx(10, 8, 7), idx(8, 10, 4), 
		idx(4, 4, 8), idx(9, 11, 12), idx(12, 10, 9), idx(10, 12, 4), idx(4, 4, 10), 
		idx(11, 13, 14), idx(14, 12, 11), idx(12, 14, 4), idx(4, 4, 12), idx(13, 15, 16), 
		idx(16, 14, 13), idx(14, 16, 4), idx(4, 4, 14), idx(15, 0, 3), idx(3, 16, 15), 
		idx(16, 3, 4), idx(4, 4, 16), idx(17, 17, 18), idx(18, 19, 17), idx(17, 17, 20), 
		idx(20, 18, 17), idx(17, 17, 21), idx(21, 20, 17), idx(17, 17, 22), idx(22, 21, 17), 
		idx(17, 17, 23), idx(23, 22, 17), idx(17, 17, 24), idx(24, 23, 17), idx(17, 17, 25), 
		idx(25, 24, 17), idx(17, 17, 19), idx(19, 25, 17)
	);

end package;
