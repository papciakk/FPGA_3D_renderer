package keyboard_inc is

	type key_t is (
		KEY_NONE,
		KEY_W,
		KEY_S,
		KEY_A,
		KEY_D,
		KEY_Q,
		KEY_E,
		KEY_Z,
		KEY_X
	);

end package keyboard_inc;
