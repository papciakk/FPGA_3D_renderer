use work.common.all;

package renderer_mesh is
	constant vertices : vertex_attr_arr_t(0 to 137) := (
		va(441, 200, 80, 11, 74, 123), va(361, 241, 102, 81, 11, 99), va(360, 243, 94, 107, 140, 2), va(440, 201, 72, 96, 148, 5), va(365, 247, 104, 156, 241, 79), va(450, 202, 80, 216, 188, 60), va(251, 237, 111, 178, 16, 90), va(250, 239, 103, 120, 140, 0), va(247, 242, 113, 75, 236, 88), va(172, 190, 102, 247, 86, 126), va(174, 193, 94, 134, 136, 0), 
		va(166, 193, 104, 20, 177, 80), va(179, 129, 80, 240, 183, 123), va(178, 131, 72, 129, 165, 6), va(170, 127, 80, 22, 98, 60), va(259, 88, 59, 171, 244, 146), va(258, 89, 51, 119, 172, 8), va(255, 82, 57, 81, 45, 40), va(369, 92, 50, 74, 239, 155), va(368, 93, 42, 105, 172, 10), va(373, 87, 48, 163, 49, 32), 
		va(445, 138, 59, 8, 168, 146), va(444, 139, 51, 97, 162, 8), va(454, 136, 57, 218, 109, 40), va(386, 255, 172, 165, 247, 111), va(491, 200, 144, 232, 187, 89), va(400, 253, 233, 172, 239, 163), va(514, 194, 202, 242, 177, 140), va(241, 249, 184, 73, 241, 121), va(243, 248, 246, 77, 234, 173), va(142, 189, 172, 10, 174, 111), 
		va(135, 182, 233, 11, 164, 163), va(147, 107, 144, 13, 84, 89), va(140, 93, 202, 14, 70, 140), va(252, 53, 115, 80, 24, 67), va(254, 34, 171, 84, 7, 117), va(396, 58, 104, 172, 30, 58), va(411, 40, 159, 180, 13, 107), va(496, 118, 115, 235, 97, 67), va(519, 105, 171, 245, 83, 117), va(397, 232, 271, 171, 205, 216), 
		va(496, 180, 244, 229, 153, 197), va(390, 215, 286, 164, 171, 239), va(476, 171, 263, 205, 134, 226), va(259, 227, 282, 92, 201, 224), va(272, 211, 296, 107, 168, 245), va(164, 170, 271, 38, 143, 216), va(191, 162, 286, 68, 126, 239), va(169, 93, 244, 40, 65, 197), va(195, 96, 263, 70, 71, 226), va(269, 41, 217, 98, 14, 178), 
		va(281, 51, 240, 111, 34, 212), va(406, 46, 206, 177, 18, 170), va(399, 55, 231, 168, 37, 206), va(501, 103, 217, 231, 76, 178), va(480, 105, 240, 207, 78, 212), va(383, 202, 291, 153, 131, 251), va(457, 164, 272, 173, 113, 244), va(337, 131, 275, 140, 97, 249), va(283, 198, 300, 125, 130, 253), va(213, 156, 291, 106, 110, 251), 
		va(217, 100, 272, 107, 83, 244), va(290, 61, 252, 127, 65, 237), va(391, 65, 244, 155, 66, 235), va(460, 107, 252, 173, 86, 237), va(165, 119, 111, 145, 98, 249), va(159, 134, 107, 71, 241, 125), va(69, 109, 110, 71, 240, 134), va(89, 98, 113, 173, 111, 244), va(41, 96, 134, 42, 220, 142), va(65, 88, 129, 241, 161, 169), 
		va(172, 125, 93, 107, 154, 4), va(67, 96, 97, 63, 131, 17), va(37, 81, 129, 10, 80, 106), va(178, 110, 97, 171, 26, 62), va(88, 85, 100, 174, 22, 72), va(60, 73, 124, 143, 8, 83), va(67, 94, 178, 63, 227, 171), va(85, 86, 166, 213, 186, 55), va(137, 104, 219, 54, 182, 215), va(140, 93, 202, 189, 180, 29), 
		va(69, 79, 181, 46, 67, 204), va(153, 92, 227, 72, 72, 227), va(86, 71, 169, 167, 8, 105), va(156, 81, 210, 141, 5, 159), va(480, 194, 160, 59, 126, 19), va(464, 214, 204, 120, 239, 186), va(542, 235, 151, 93, 246, 156), va(540, 216, 129, 35, 113, 39), va(582, 249, 85, 73, 240, 110), va(562, 232, 80, 31, 114, 44), 
		va(489, 182, 227, 212, 139, 219), va(572, 219, 158, 225, 147, 205), va(618, 247, 80, 214, 134, 218), va(505, 162, 182, 217, 37, 125), va(570, 200, 136, 199, 27, 93), va(598, 230, 76, 177, 33, 57), va(595, 252, 78, 112, 227, 50), va(573, 236, 76, 114, 166, 7), va(586, 246, 83, 213, 37, 101), va(572, 235, 80, 236, 163, 180), 
		va(630, 252, 74, 234, 182, 89), va(609, 245, 80, 76, 137, 10), va(608, 236, 72, 188, 104, 18), va(595, 234, 78, 119, 245, 172), va(302, 175, 20, 113, 156, 4), va(315, 190, 38, 165, 247, 114), va(334, 181, 33, 233, 186, 91), va(314, 180, 59, 157, 241, 80), va(325, 174, 56, 216, 188, 61), va(290, 189, 40, 73, 242, 123), 
		va(298, 179, 60, 75, 236, 88), va(272, 179, 38, 9, 174, 114), va(287, 172, 59, 20, 177, 80), va(273, 164, 33, 12, 84, 91), va(288, 164, 56, 22, 97, 61), va(292, 155, 28, 80, 23, 69), va(299, 158, 53, 81, 44, 41), va(317, 156, 26, 172, 29, 60), va(315, 158, 52, 163, 49, 33), va(335, 166, 28, 236, 96, 69), 
		va(326, 165, 53, 218, 108, 41), va(339, 212, 81, 125, 187, 15), va(385, 187, 68, 145, 170, 9), va(358, 236, 101, 127, 190, 16), va(432, 197, 80, 148, 171, 10), va(274, 209, 86, 99, 186, 18), va(255, 232, 109, 98, 188, 19), va(229, 182, 81, 81, 166, 15), va(185, 189, 101, 78, 167, 16), va(231, 146, 68, 81, 140, 9), 
		va(189, 132, 80, 79, 139, 10), va(278, 121, 56, 101, 123, 2), va(263, 93, 60, 100, 120, 3), va(343, 124, 50, 127, 125, 0), va(365, 97, 52, 129, 121, 0), va(388, 151, 56, 146, 144, 2), va(435, 140, 60, 149, 143, 3)
	);

	constant indices : indices_arr_t(0 to 255) := (
		idx(0, 1, 2), idx(2, 3, 0), 
		idx(3, 2, 4), idx(4, 5, 3), idx(1, 6, 7), idx(7, 2, 1), idx(2, 7, 8), idx(8, 4, 2), idx(6, 9, 10), idx(10, 7, 6), idx(7, 10, 11), idx(11, 8, 7), 
		idx(9, 12, 13), idx(13, 10, 9), idx(10, 13, 14), idx(14, 11, 10), idx(12, 15, 16), idx(16, 13, 12), idx(13, 16, 17), idx(17, 14, 13), idx(15, 18, 19), idx(19, 16, 15), 
		idx(16, 19, 20), idx(20, 17, 16), idx(18, 21, 22), idx(22, 19, 18), idx(19, 22, 23), idx(23, 20, 19), idx(21, 0, 3), idx(3, 22, 21), idx(22, 3, 5), idx(5, 23, 22), 
		idx(5, 4, 24), idx(24, 25, 5), idx(25, 24, 26), idx(26, 27, 25), idx(4, 8, 28), idx(28, 24, 4), idx(24, 28, 29), idx(29, 26, 24), idx(8, 11, 30), idx(30, 28, 8), 
		idx(28, 30, 31), idx(31, 29, 28), idx(11, 14, 32), idx(32, 30, 11), idx(30, 32, 33), idx(33, 31, 30), idx(14, 17, 34), idx(34, 32, 14), idx(32, 34, 35), idx(35, 33, 32), 
		idx(17, 20, 36), idx(36, 34, 17), idx(34, 36, 37), idx(37, 35, 34), idx(20, 23, 38), idx(38, 36, 20), idx(36, 38, 39), idx(39, 37, 36), idx(23, 5, 25), idx(25, 38, 23), 
		idx(38, 25, 27), idx(27, 39, 38), idx(27, 26, 40), idx(40, 41, 27), idx(41, 40, 42), idx(42, 43, 41), idx(26, 29, 44), idx(44, 40, 26), idx(40, 44, 45), idx(45, 42, 40), 
		idx(29, 31, 46), idx(46, 44, 29), idx(44, 46, 47), idx(47, 45, 44), idx(31, 33, 48), idx(48, 46, 31), idx(46, 48, 49), idx(49, 47, 46), idx(33, 35, 50), idx(50, 48, 33), 
		idx(48, 50, 51), idx(51, 49, 48), idx(35, 37, 52), idx(52, 50, 35), idx(50, 52, 53), idx(53, 51, 50), idx(37, 39, 54), idx(54, 52, 37), idx(52, 54, 55), idx(55, 53, 52), 
		idx(39, 27, 41), idx(41, 54, 39), idx(54, 41, 43), idx(43, 55, 54), idx(43, 42, 56), idx(56, 57, 43), idx(57, 56, 58), idx(58, 58, 57), idx(42, 45, 59), idx(59, 56, 42), 
		idx(56, 59, 58), idx(58, 58, 56), idx(45, 47, 60), idx(60, 59, 45), idx(59, 60, 58), idx(58, 58, 59), idx(47, 49, 61), idx(61, 60, 47), idx(60, 61, 58), idx(58, 58, 60), 
		idx(49, 51, 62), idx(62, 61, 49), idx(61, 62, 58), idx(58, 58, 61), idx(51, 53, 63), idx(63, 62, 51), idx(62, 63, 58), idx(58, 58, 62), idx(53, 55, 64), idx(64, 63, 53), 
		idx(63, 64, 58), idx(58, 58, 63), idx(55, 43, 57), idx(57, 64, 55), idx(64, 57, 58), idx(58, 58, 64), idx(65, 66, 67), idx(67, 68, 65), idx(68, 67, 69), idx(69, 70, 68), 
		idx(66, 71, 72), idx(72, 67, 66), idx(67, 72, 73), idx(73, 69, 67), idx(71, 74, 75), idx(75, 72, 71), idx(72, 75, 76), idx(76, 73, 72), idx(74, 65, 68), idx(68, 75, 74), 
		idx(75, 68, 70), idx(70, 76, 75), idx(70, 69, 77), idx(77, 78, 70), idx(78, 77, 79), idx(79, 80, 78), idx(69, 73, 81), idx(81, 77, 69), idx(77, 81, 82), idx(82, 79, 77), 
		idx(73, 76, 83), idx(83, 81, 73), idx(81, 83, 84), idx(84, 82, 81), idx(76, 70, 78), idx(78, 83, 76), idx(83, 78, 80), idx(80, 84, 83), idx(85, 86, 87), idx(87, 88, 85), 
		idx(88, 87, 89), idx(89, 90, 88), idx(86, 91, 92), idx(92, 87, 86), idx(87, 92, 93), idx(93, 89, 87), idx(91, 94, 95), idx(95, 92, 91), idx(92, 95, 96), idx(96, 93, 92), 
		idx(94, 85, 88), idx(88, 95, 94), idx(95, 88, 90), idx(90, 96, 95), idx(90, 89, 97), idx(97, 98, 90), idx(98, 97, 99), idx(99, 100, 98), idx(89, 93, 101), idx(101, 97, 89), 
		idx(97, 101, 102), idx(102, 99, 97), idx(93, 96, 103), idx(103, 101, 93), idx(101, 103, 104), idx(104, 102, 101), idx(96, 90, 98), idx(98, 103, 96), idx(103, 98, 100), idx(100, 104, 103), 
		idx(105, 105, 106), idx(106, 107, 105), idx(107, 106, 108), idx(108, 109, 107), idx(105, 105, 110), idx(110, 106, 105), idx(106, 110, 111), idx(111, 108, 106), idx(105, 105, 112), idx(112, 110, 105), 
		idx(110, 112, 113), idx(113, 111, 110), idx(105, 105, 114), idx(114, 112, 105), idx(112, 114, 115), idx(115, 113, 112), idx(105, 105, 116), idx(116, 114, 105), idx(114, 116, 117), idx(117, 115, 114), 
		idx(105, 105, 118), idx(118, 116, 105), idx(116, 118, 119), idx(119, 117, 116), idx(105, 105, 120), idx(120, 118, 105), idx(118, 120, 121), idx(121, 119, 118), idx(105, 105, 107), idx(107, 120, 105), 
		idx(120, 107, 109), idx(109, 121, 120), idx(109, 108, 122), idx(122, 123, 109), idx(123, 122, 124), idx(124, 125, 123), idx(108, 111, 126), idx(126, 122, 108), idx(122, 126, 127), idx(127, 124, 122), 
		idx(111, 113, 128), idx(128, 126, 111), idx(126, 128, 129), idx(129, 127, 126), idx(113, 115, 130), idx(130, 128, 113), idx(128, 130, 131), idx(131, 129, 128), idx(115, 117, 132), idx(132, 130, 115), 
		idx(130, 132, 133), idx(133, 131, 130), idx(117, 119, 134), idx(134, 132, 117), idx(132, 134, 135), idx(135, 133, 132), idx(119, 121, 136), idx(136, 134, 119), idx(134, 136, 137), idx(137, 135, 134), 
		idx(121, 109, 123), idx(123, 136, 121), idx(136, 123, 125), idx(125, 137, 136)
	);

end package renderer_mesh;
