use work.definitions.all;

package mesh is
	constant vertices : vertex_attr_arr_t(0 to 85) := (
		va(-14, 0, 22936, 0, 0, 32767), va(-14, 9954, 20664, 0, 15038, 29112), va(-4333, 8969, 20664, -6525, 13549, 29112), 
		va(-7797, 6206, 20664, -11757, 9376, 29112), va(-9719, 2215, 20664, -14661, 3346, 29112), va(-9719, -2215, 20664, -14661, -3346, 29112), 
		va(-7797, -6206, 20664, -11757, -9376, 29112), va(-4333, -8969, 20664, -6525, -13549, 29112), va(-14, -9954, 20664, 0, -15038, 29112), 
		va(4304, -8969, 20664, 6525, -13549, 29112), va(7768, -6206, 20664, 11757, -9376, 29112), va(9690, -2215, 20664, 14661, -3346, 29112), 
		va(9690, 2215, 20664, 14661, 3346, 29112), va(7768, 6206, 20664, 11757, 9376, 29112), va(4304, 8969, 20664, 6525, 13549, 29112), 
		va(-14, 17938, 14297, 0, 26002, 19939), va(-7797, 16161, 14297, -11282, 23427, 19939), va(-14039, 11184, 14297, -20329, 16212, 19939), 
		va(-17502, 3991, 14297, -25350, 5786, 19939), va(-17502, -3991, 14297, -25350, -5786, 19939), va(-14039, -11184, 14297, -20329, -16212, 19939), 
		va(-7797, -16161, 14297, -11282, -23427, 19939), va(-14, -17938, 14297, 0, -26002, 19939), va(7768, -16161, 14297, 11282, -23427, 19939), 
		va(14010, -11184, 14297, 20329, -16212, 19939), va(17473, -3991, 14297, 25350, -5786, 19939), va(17473, 3991, 14297, 25350, 5786, 19939), 
		va(14010, 11184, 14297, 20329, 16212, 19939), va(7768, 16161, 14297, 11282, 23427, 19939), va(-14, 22368, 5097, 0, 31994, 7077), 
		va(-9719, 20153, 5097, -13882, 28825, 7077), va(-17502, 13946, 5097, -25014, 19948, 7077), va(-21822, 4977, 5097, -31192, 7119, 7077), 
		va(-21822, -4977, 5097, -31192, -7119, 7077), va(-17502, -13946, 5097, -25014, -19948, 7077), va(-9719, -20153, 5097, -13882, -28825, 7077), 
		va(-14, -22368, 5097, 0, -31994, 7077), va(9690, -20153, 5097, 13882, -28825, 7077), va(17473, -13946, 5097, 25014, -19948, 7077), 
		va(21793, -4977, 5097, 31192, -7119, 7077), va(21793, 4977, 5097, 31192, 7119, 7077), va(17473, 13946, 5097, 25014, 19948, 7077), 
		va(9690, 20153, 5097, 13882, 28825, 7077), va(-14, 22368, -5112, 0, 31994, -7077), va(-9719, 20153, -5112, -13882, 28825, -7077), 
		va(-17502, 13946, -5112, -25014, 19948, -7077), va(-21822, 4977, -5112, -31192, 7119, -7077), va(-21822, -4977, -5112, -31192, -7119, -7077), 
		va(-17502, -13946, -5112, -25014, -19948, -7077), va(-9719, -20153, -5112, -13882, -28825, -7077), va(-14, -22368, -5112, 0, -31994, -7077), 
		va(9690, -20153, -5112, 13882, -28825, -7077), va(17473, -13946, -5112, 25014, -19948, -7077), va(21793, -4977, -5112, 31192, -7119, -7077), 
		va(21793, 4977, -5112, 31192, 7119, -7077), va(17473, 13946, -5112, 25014, 19948, -7077), va(9690, 20153, -5112, 13882, 28825, -7077), 
		va(-14, 17938, -14312, 0, 26002, -19939), va(-7797, 16161, -14312, -11282, 23427, -19939), va(-14039, 11184, -14312, -20329, 16212, -19939), 
		va(-17502, 3991, -14312, -25350, 5786, -19939), va(-17502, -3991, -14312, -25350, -5786, -19939), va(-14039, -11184, -14312, -20329, -16212, -19939), 
		va(-7797, -16161, -14312, -11282, -23427, -19939), va(-14, -17938, -14312, 0, -26002, -19939), va(7768, -16161, -14312, 11282, -23427, -19939), 
		va(14010, -11184, -14312, 20329, -16212, -19939), va(17473, -3991, -14312, 25350, -5786, -19939), va(17473, 3991, -14312, 25350, 5786, -19939), 
		va(14010, 11184, -14312, 20329, 16212, -19939), va(7768, 16161, -14312, 11282, 23427, -19939), va(-14, 9954, -20679, 0, 15038, -29112), 
		va(-4333, 8969, -20679, -6525, 13549, -29112), va(-7797, 6206, -20679, -11757, 9376, -29112), va(-9719, 2215, -20679, -14661, 3346, -29112), 
		va(-9719, -2215, -20679, -14661, -3346, -29112), va(-7797, -6206, -20679, -11757, -9376, -29112), va(-4333, -8969, -20679, -6525, -13549, -29112), 
		va(-14, -9954, -20679, 0, -15038, -29112), va(4304, -8969, -20679, 6525, -13549, -29112), va(7768, -6206, -20679, 11757, -9376, -29112), 
		va(9690, -2215, -20679, 14661, -3346, -29112), va(9690, 2215, -20679, 14661, 3346, -29112), va(7768, 6206, -20679, 11757, 9376, -29112), 
		va(4304, 8969, -20679, 6525, 13549, -29112), va(-14, 0, -22951, 0, 0, -32767)
	);

	constant indices : indices_arr_t(0 to 167) := (
		idx(0, 1, 2), idx(0, 2, 3), idx(0, 3, 4), idx(0, 4, 5), idx(0, 5, 6), 
		idx(0, 6, 7), idx(0, 7, 8), idx(0, 8, 9), idx(0, 9, 10), idx(0, 10, 11), 
		idx(0, 11, 12), idx(0, 12, 13), idx(0, 13, 14), idx(0, 14, 1), idx(1, 15, 16), 
		idx(1, 16, 2), idx(2, 16, 17), idx(2, 17, 3), idx(3, 17, 18), idx(3, 18, 4), 
		idx(4, 18, 19), idx(4, 19, 5), idx(5, 19, 20), idx(5, 20, 6), idx(6, 20, 21), 
		idx(6, 21, 7), idx(7, 21, 22), idx(7, 22, 8), idx(8, 22, 23), idx(8, 23, 9), 
		idx(9, 23, 24), idx(9, 24, 10), idx(10, 24, 25), idx(10, 25, 11), idx(11, 25, 26), 
		idx(11, 26, 12), idx(12, 26, 27), idx(12, 27, 13), idx(13, 27, 28), idx(13, 28, 14), 
		idx(14, 28, 15), idx(14, 15, 1), idx(15, 29, 30), idx(15, 30, 16), idx(16, 30, 31), 
		idx(16, 31, 17), idx(17, 31, 32), idx(17, 32, 18), idx(18, 32, 33), idx(18, 33, 19), 
		idx(19, 33, 34), idx(19, 34, 20), idx(20, 34, 35), idx(20, 35, 21), idx(21, 35, 36), 
		idx(21, 36, 22), idx(22, 36, 37), idx(22, 37, 23), idx(23, 37, 38), idx(23, 38, 24), 
		idx(24, 38, 39), idx(24, 39, 25), idx(25, 39, 40), idx(25, 40, 26), idx(26, 40, 41), 
		idx(26, 41, 27), idx(27, 41, 42), idx(27, 42, 28), idx(28, 42, 29), idx(28, 29, 15), 
		idx(29, 43, 44), idx(29, 44, 30), idx(30, 44, 45), idx(30, 45, 31), idx(31, 45, 46), 
		idx(31, 46, 32), idx(32, 46, 47), idx(32, 47, 33), idx(33, 47, 48), idx(33, 48, 34), 
		idx(34, 48, 49), idx(34, 49, 35), idx(35, 49, 50), idx(35, 50, 36), idx(36, 50, 51), 
		idx(36, 51, 37), idx(37, 51, 52), idx(37, 52, 38), idx(38, 52, 53), idx(38, 53, 39), 
		idx(39, 53, 54), idx(39, 54, 40), idx(40, 54, 55), idx(40, 55, 41), idx(41, 55, 56), 
		idx(41, 56, 42), idx(42, 56, 43), idx(42, 43, 29), idx(43, 57, 58), idx(43, 58, 44), 
		idx(44, 58, 59), idx(44, 59, 45), idx(45, 59, 60), idx(45, 60, 46), idx(46, 60, 61), 
		idx(46, 61, 47), idx(47, 61, 62), idx(47, 62, 48), idx(48, 62, 63), idx(48, 63, 49), 
		idx(49, 63, 64), idx(49, 64, 50), idx(50, 64, 65), idx(50, 65, 51), idx(51, 65, 66), 
		idx(51, 66, 52), idx(52, 66, 67), idx(52, 67, 53), idx(53, 67, 68), idx(53, 68, 54), 
		idx(54, 68, 69), idx(54, 69, 55), idx(55, 69, 70), idx(55, 70, 56), idx(56, 70, 57), 
		idx(56, 57, 43), idx(57, 71, 72), idx(57, 72, 58), idx(58, 72, 73), idx(58, 73, 59), 
		idx(59, 73, 74), idx(59, 74, 60), idx(60, 74, 75), idx(60, 75, 61), idx(61, 75, 76), 
		idx(61, 76, 62), idx(62, 76, 77), idx(62, 77, 63), idx(63, 77, 78), idx(63, 78, 64), 
		idx(64, 78, 79), idx(64, 79, 65), idx(65, 79, 80), idx(65, 80, 66), idx(66, 80, 81), 
		idx(66, 81, 67), idx(67, 81, 82), idx(67, 82, 68), idx(68, 82, 83), idx(68, 83, 69), 
		idx(69, 83, 84), idx(69, 84, 70), idx(70, 84, 71), idx(70, 71, 57), idx(85, 72, 71), 
		idx(85, 73, 72), idx(85, 74, 73), idx(85, 75, 74), idx(85, 76, 75), idx(85, 77, 76), 
		idx(85, 78, 77), idx(85, 79, 78), idx(85, 80, 79), idx(85, 81, 80), idx(85, 82, 81), 
		idx(85, 83, 82), idx(85, 84, 83), idx(85, 71, 84)
	);

end package;
