use work.definitions.all;

package mesh is
	constant vertices : vertex_attr_arr_t(0 to 137) := (
		va(8463, 5887, -19, -32751, 1040, 0), va(5565, 5887, 7073, -23158, 1044, -23158), va(5581, 6589, 7089, -3165, 32460, -3165), 
		va(8485, 6589, -19, -4641, 32437, 0), va(6072, 5887, 7580, 19449, 17808, 19449), va(9176, 5887, -19, 27525, 17777, 0), 
		va(-1527, 5887, 9970, -34, 927, -32754), va(-1527, 6589, 9993, -25, 32435, -4655), va(-1527, 5887, 10684, 0, 17777, 27525), 
		va(-8861, 5887, 7073, 23816, -5808, -21743), va(-8666, 6589, 7089, 2673, 31878, -7095), va(-9127, 5887, 7580, -19492, 17634, 19565), 
		va(-11518, 5887, -19, 32747, 1040, 486), va(-11540, 6589, -19, 4903, 32395, 441), va(-12231, 5887, -19, -27533, 17766, -15), 
		va(-8620, 5887, -7113, 23158, 1044, 23158), va(-8636, 6589, -7129, 3165, 32460, 3165), va(-9127, 5887, -7619, -19449, 17808, -19449), 
		va(-1527, 5887, -10010, 0, 1040, 32751), va(-1527, 6589, -10032, 0, 32437, 4641), va(-1527, 5887, -10724, 0, 17777, -27525), 
		va(5565, 5887, -7113, -23158, 1044, 23158), va(5581, 6589, -7129, -3165, 32460, 3165), va(6072, 5887, -7619, 19449, 17808, -19449), 
		va(7814, 334, 9321, 22078, 9940, 22078), va(11629, 334, -19, 31232, 9911, 0), va(8605, -4816, 10113, 23027, -3627, 23027), 
		va(12744, -4816, -19, 32566, -3622, 0), va(-1527, 334, 13137, 0, 9911, 31232), va(-1527, -4816, 14252, 0, -3622, 32566), 
		va(-10869, 334, 9321, -22078, 9940, 22078), va(-11661, -4816, 10113, -23027, -3627, 23027), va(-14684, 334, -19, -31232, 9911, 0), 
		va(-15799, -4816, -19, -32566, -3622, 0), va(-10869, 334, -9361, -22078, 9940, -22078), va(-11661, -4816, -10153, -23027, -3627, -23027), 
		va(-1527, 334, -13177, 0, 9911, -31232), va(-1527, -4816, -14292, 0, -3622, -32566), va(7814, 334, -9361, 22078, 9940, -22078), 
		va(8605, -4816, -10153, 23027, -3627, -23027), va(7339, -8496, 8846, 18980, -18793, 18980), va(10960, -8496, -19, 26864, -18762, 0), 
		va(6072, -10169, 7580, 13622, -26506, 13622), va(9176, -10169, -19, 19293, -26485, 0), va(-1527, -8496, 12468, 0, -18762, 26864), 
		va(-1527, -10169, 10684, 0, -26485, 19293), va(-10394, -8496, 8846, -18980, -18793, 18980), va(-9127, -10169, 7580, -13622, -26506, 13622), 
		va(-14015, -8496, -19, -26864, -18762, 0), va(-12231, -10169, -19, -19293, -26485, 0), va(-10394, -8496, -8886, -18980, -18793, -18980), 
		va(-9127, -10169, -7619, -13622, -26506, -13622), va(-1527, -8496, -12508, 0, -18762, -26864), va(-1527, -10169, -10724, 0, -26485, -19293), 
		va(7339, -8496, -8886, 18980, -18793, -18980), va(6072, -10169, -7619, 13622, -26506, -13622), va(4979, -10905, 6487, 6607, -31406, 6607), 
		va(7637, -10905, -19, 9339, -31408, 0), va(-1527, -11239, -19, 0, -32767, 0), va(-1527, -10905, 9145, 0, -31408, 9339), 
		va(-8035, -10905, 6487, -6607, -31406, 6607), va(-10693, -10905, -19, -9339, -31408, 0), va(-8035, -10905, -6527, -6607, -31406, -6607), 
		va(-1527, -10905, -9185, 0, -31408, -9339), va(4979, -10905, -6527, 6607, -31406, -6607), va(-12945, 3211, -19, 1258, -32743, -100), 
		va(-12588, 4014, 1585, -596, 8936, 31519), va(-19501, 3713, 1585, -622, 6707, 32067), va(-18743, 3010, -19, 9230, -31437, -474), 
		va(-21865, 1605, 1585, -9628, 4143, 31045), va(-20795, 1605, -19, 30551, -11765, -1382), va(-12231, 4816, -19, -1550, 32730, 48), 
		va(-20260, 4415, -19, -14485, 29389, 415), va(-22936, 1605, -19, -32306, 5467, 347), va(-12588, 4014, -1625, -581, 8799, -31558), 
		va(-19501, 3713, -1625, -318, 5852, -32239), va(-21865, 1605, -1625, -8961, 3320, -31342), va(-20327, -2291, 1585, -3987, -3269, 32359), 
		va(-19635, -1605, -19, 26792, 18859, -453), va(-15443, -5887, 1585, -10984, -16585, 26038), va(-15799, -4816, -19, 20367, 25650, -965), 
		va(-21018, -2977, -19, -25385, -20717, 258), va(-15086, -6957, -19, -18714, -26896, 249), va(-20327, -2291, -1625, -3458, -2913, -32454), 
		va(-15443, -5887, -1625, -9860, -15953, -26870), va(10603, -1070, -19, -15931, 28633, -241), va(10603, -4014, 3512, 10718, -7805, 29965), 
		va(16580, 334, 2415, 5226, 805, 32338), va(15510, 1605, -19, -22837, 23485, 774), va(19881, 5887, 1318, -205, 12492, 30292), 
		va(17740, 5887, -19, -23704, 22548, 1843), va(10603, -6957, -19, 21422, -24795, -81), va(17650, -936, -19, 25156, -20989, -566), 
		va(22021, 5887, -19, 21184, -24955, -1465), va(10603, -4014, -3552, 11324, -7679, -29774), va(16580, 334, -2455, 6047, 266, -32203), 
		va(19881, 5887, -1357, 1657, 10336, -31050), va(20784, 6364, 1050, 7598, 25537, 19074), va(18632, 6288, -19, 1361, 32657, 2308), 
		va(19881, 5887, 782, 10348, -1488, -31054), va(18453, 5887, -19, 29526, -14201, 443), va(22936, 6439, -19, 31237, 9821, -1217), 
		va(21308, 5887, -19, -10546, 31023, -106), va(20784, 6364, -1090, 11978, 23899, -18949), va(19881, 5887, -822, 11121, -3846, 30581), 
		va(-1527, 11239, -19, 0, 32767, 0), va(121, 10035, 1628, 22197, 9406, 22192), va(791, 10035, -19, 31376, 9445, 4), 
		va(-514, 8028, 993, 19513, 17681, 19502), va(-100, 8028, -19, 27642, 17596, 8), va(-1527, 10035, 2299, -4, 9445, 31376), 
		va(-1527, 8028, 1407, -8, 17596, 27642), va(-3176, 10035, 1628, -22192, 9406, 22197), va(-2540, 8028, 993, -19502, 17681, 19513), 
		va(-3846, 10035, -19, -31376, 9445, -4), va(-2954, 8028, -19, -27642, 17596, -8), va(-3176, 10035, -1668, -22197, 9406, -22192), 
		va(-2540, 8028, -1033, -19513, 17681, -19502), va(-1527, 10035, -2339, 4, 9445, -31376), va(-1527, 8028, -1447, 8, 17596, -27642), 
		va(121, 10035, -1668, 22192, 9406, -22197), va(-514, 8028, -1033, 19502, 17681, -19513), va(2652, 6957, 4160, 6362, 31507, 6362), 
		va(4359, 6957, -19, 9025, 31500, 0), va(5059, 5887, 6566, 6951, 31258, 6951), va(7749, 5887, -19, 9867, 31246, 0), 
		va(-1527, 6957, 5867, 0, 31500, 9025), va(-1527, 5887, 9257, 0, 31246, 9867), va(-5707, 6957, 4160, -6362, 31507, 6362), 
		va(-8114, 5887, 6566, -6951, 31258, 6951), va(-7414, 6957, -19, -9025, 31500, 0), va(-10804, 5887, -19, -9867, 31246, 0), 
		va(-5707, 6957, -4199, -6362, 31507, -6362), va(-8114, 5887, -6606, -6951, 31258, -6951), va(-1527, 6957, -5907, 0, 31500, -9025), 
		va(-1527, 5887, -9296, 0, 31246, -9867), va(2652, 6957, -4199, 6362, 31507, -6362), va(5059, 5887, -6606, 6951, 31258, -6951)
		
	);

	constant indices : indices_arr_t(0 to 255) := (
		idx(0, 1, 2), idx(2, 3, 0), idx(3, 2, 4), idx(4, 5, 3), idx(1, 6, 7), 
		idx(7, 2, 1), idx(2, 7, 8), idx(8, 4, 2), idx(6, 9, 10), idx(10, 7, 6), 
		idx(7, 10, 11), idx(11, 8, 7), idx(9, 12, 13), idx(13, 10, 9), idx(10, 13, 14), 
		idx(14, 11, 10), idx(12, 15, 16), idx(16, 13, 12), idx(13, 16, 17), idx(17, 14, 13), 
		idx(15, 18, 19), idx(19, 16, 15), idx(16, 19, 20), idx(20, 17, 16), idx(18, 21, 22), 
		idx(22, 19, 18), idx(19, 22, 23), idx(23, 20, 19), idx(21, 0, 3), idx(3, 22, 21), 
		idx(22, 3, 5), idx(5, 23, 22), idx(5, 4, 24), idx(24, 25, 5), idx(25, 24, 26), 
		idx(26, 27, 25), idx(4, 8, 28), idx(28, 24, 4), idx(24, 28, 29), idx(29, 26, 24), 
		idx(8, 11, 30), idx(30, 28, 8), idx(28, 30, 31), idx(31, 29, 28), idx(11, 14, 32), 
		idx(32, 30, 11), idx(30, 32, 33), idx(33, 31, 30), idx(14, 17, 34), idx(34, 32, 14), 
		idx(32, 34, 35), idx(35, 33, 32), idx(17, 20, 36), idx(36, 34, 17), idx(34, 36, 37), 
		idx(37, 35, 34), idx(20, 23, 38), idx(38, 36, 20), idx(36, 38, 39), idx(39, 37, 36), 
		idx(23, 5, 25), idx(25, 38, 23), idx(38, 25, 27), idx(27, 39, 38), idx(27, 26, 40), 
		idx(40, 41, 27), idx(41, 40, 42), idx(42, 43, 41), idx(26, 29, 44), idx(44, 40, 26), 
		idx(40, 44, 45), idx(45, 42, 40), idx(29, 31, 46), idx(46, 44, 29), idx(44, 46, 47), 
		idx(47, 45, 44), idx(31, 33, 48), idx(48, 46, 31), idx(46, 48, 49), idx(49, 47, 46), 
		idx(33, 35, 50), idx(50, 48, 33), idx(48, 50, 51), idx(51, 49, 48), idx(35, 37, 52), 
		idx(52, 50, 35), idx(50, 52, 53), idx(53, 51, 50), idx(37, 39, 54), idx(54, 52, 37), 
		idx(52, 54, 55), idx(55, 53, 52), idx(39, 27, 41), idx(41, 54, 39), idx(54, 41, 43), 
		idx(43, 55, 54), idx(43, 42, 56), idx(56, 57, 43), idx(57, 56, 58), idx(58, 58, 57), 
		idx(42, 45, 59), idx(59, 56, 42), idx(56, 59, 58), idx(58, 58, 56), idx(45, 47, 60), 
		idx(60, 59, 45), idx(59, 60, 58), idx(58, 58, 59), idx(47, 49, 61), idx(61, 60, 47), 
		idx(60, 61, 58), idx(58, 58, 60), idx(49, 51, 62), idx(62, 61, 49), idx(61, 62, 58), 
		idx(58, 58, 61), idx(51, 53, 63), idx(63, 62, 51), idx(62, 63, 58), idx(58, 58, 62), 
		idx(53, 55, 64), idx(64, 63, 53), idx(63, 64, 58), idx(58, 58, 63), idx(55, 43, 57), 
		idx(57, 64, 55), idx(64, 57, 58), idx(58, 58, 64), idx(65, 66, 67), idx(67, 68, 65), 
		idx(68, 67, 69), idx(69, 70, 68), idx(66, 71, 72), idx(72, 67, 66), idx(67, 72, 73), 
		idx(73, 69, 67), idx(71, 74, 75), idx(75, 72, 71), idx(72, 75, 76), idx(76, 73, 72), 
		idx(74, 65, 68), idx(68, 75, 74), idx(75, 68, 70), idx(70, 76, 75), idx(70, 69, 77), 
		idx(77, 78, 70), idx(78, 77, 79), idx(79, 80, 78), idx(69, 73, 81), idx(81, 77, 69), 
		idx(77, 81, 82), idx(82, 79, 77), idx(73, 76, 83), idx(83, 81, 73), idx(81, 83, 84), 
		idx(84, 82, 81), idx(76, 70, 78), idx(78, 83, 76), idx(83, 78, 80), idx(80, 84, 83), 
		idx(85, 86, 87), idx(87, 88, 85), idx(88, 87, 89), idx(89, 90, 88), idx(86, 91, 92), 
		idx(92, 87, 86), idx(87, 92, 93), idx(93, 89, 87), idx(91, 94, 95), idx(95, 92, 91), 
		idx(92, 95, 96), idx(96, 93, 92), idx(94, 85, 88), idx(88, 95, 94), idx(95, 88, 90), 
		idx(90, 96, 95), idx(90, 89, 97), idx(97, 98, 90), idx(98, 97, 99), idx(99, 100, 98), 
		idx(89, 93, 101), idx(101, 97, 89), idx(97, 101, 102), idx(102, 99, 97), idx(93, 96, 103), 
		idx(103, 101, 93), idx(101, 103, 104), idx(104, 102, 101), idx(96, 90, 98), idx(98, 103, 96), 
		idx(103, 98, 100), idx(100, 104, 103), idx(105, 105, 106), idx(106, 107, 105), idx(107, 106, 108), 
		idx(108, 109, 107), idx(105, 105, 110), idx(110, 106, 105), idx(106, 110, 111), idx(111, 108, 106), 
		idx(105, 105, 112), idx(112, 110, 105), idx(110, 112, 113), idx(113, 111, 110), idx(105, 105, 114), 
		idx(114, 112, 105), idx(112, 114, 115), idx(115, 113, 112), idx(105, 105, 116), idx(116, 114, 105), 
		idx(114, 116, 117), idx(117, 115, 114), idx(105, 105, 118), idx(118, 116, 105), idx(116, 118, 119), 
		idx(119, 117, 116), idx(105, 105, 120), idx(120, 118, 105), idx(118, 120, 121), idx(121, 119, 118), 
		idx(105, 105, 107), idx(107, 120, 105), idx(120, 107, 109), idx(109, 121, 120), idx(109, 108, 122), 
		idx(122, 123, 109), idx(123, 122, 124), idx(124, 125, 123), idx(108, 111, 126), idx(126, 122, 108), 
		idx(122, 126, 127), idx(127, 124, 122), idx(111, 113, 128), idx(128, 126, 111), idx(126, 128, 129), 
		idx(129, 127, 126), idx(113, 115, 130), idx(130, 128, 113), idx(128, 130, 131), idx(131, 129, 128), 
		idx(115, 117, 132), idx(132, 130, 115), idx(130, 132, 133), idx(133, 131, 130), idx(117, 119, 134), 
		idx(134, 132, 117), idx(132, 134, 135), idx(135, 133, 132), idx(119, 121, 136), idx(136, 134, 119), 
		idx(134, 136, 137), idx(137, 135, 134), idx(121, 109, 123), idx(123, 136, 121), idx(136, 123, 125), 
		idx(125, 137, 136)
	);

end package;
