use work.common.all;

package renderer_mesh is
	constant vertices : vertex_attr_arr_t(0 to 301) := (
		va(9326, 7693, -3126, 1, 108, 139), va(7910, 10609, 1355, 18, 74, 86), va(7807, 11127, 945, 49, 178, 40), va(9205, 8247, -3482, 37, 202, 77), va(8121, 11229, 1102, 181, 236, 93), va(9567, 8247, -3482, 190, 219, 66), va(8561, 10814, 1674, 221, 211, 137), va(10073, 7693, -3126, 236, 181, 91), va(4150, 12657, 4506, 64, 49, 48), va(4096, 13151, 4060, 82, 160, 12), va(4277, 13326, 4325, 158, 249, 112), 
		va(4536, 13013, 5048, 181, 232, 170), va(-1192, 13434, 5693, 126, 39, 34), va(-1192, 13922, 5235, 126, 153, 2), va(-1192, 14121, 5542, 127, 253, 119), va(-1192, 13844, 6325, 127, 240, 183), va(-6837, 12669, 4506, 190, 36, 64), va(-6566, 13163, 4060, 170, 151, 10), va(-6669, 13332, 4325, 95, 249, 112), va(-6916, 13019, 5048, 72, 232, 171), va(-10446, 10621, 1355, 233, 63, 99), 
		va(-10235, 11139, 945, 209, 171, 41), va(-10512, 11241, 1102, 72, 236, 93), va(-10946, 10832, 1674, 32, 211, 137), va(-11717, 7711, -3126, 251, 108, 140), va(-11597, 8259, -3482, 216, 202, 79), va(-11958, 8259, -3482, 64, 219, 66), va(-12464, 7711, -3126, 17, 181, 91), va(-10302, 4795, -7609, 235, 142, 191), va(-10193, 5380, -7916, 204, 226, 115), va(-10506, 5277, -8066, 72, 202, 40), 
		va(-10946, 4590, -7928, 32, 151, 45), va(-6542, 2747, -10753, 189, 167, 230), va(-6482, 3355, -11031, 171, 244, 142), va(-6669, 3181, -11290, 95, 189, 21), va(-6928, 2391, -11302, 72, 129, 12), va(-1198, 1970, -11946, 127, 176, 244), va(-1198, 2584, -12205, 127, 251, 152), va(-1198, 2385, -12507, 127, 185, 14), va(-1198, 1560, -12573, 127, 121, 0), va(4144, 2735, -10753, 64, 167, 230), 
		va(4084, 3343, -11031, 82, 244, 142), va(4271, 3174, -11290, 158, 189, 21), va(4530, 2385, -11302, 181, 129, 12), va(7904, 4783, -7609, 18, 142, 191), va(7801, 5367, -7916, 49, 227, 115), va(8115, 5265, -8066, 181, 202, 40), va(8554, 4572, -7928, 221, 151, 45), va(10121, 8024, 4584, 228, 199, 149), va(11880, 4404, -988, 244, 167, 100), va(11320, 5229, 7247, 233, 186, 161), 
		va(13272, 1216, 1084, 250, 153, 109), va(11802, 2403, 9422, 236, 152, 185), va(13826, -1759, 3018, 253, 117, 132), va(5452, 10573, 8500, 185, 222, 186), va(6157, 8048, 11579, 188, 211, 199), va(6440, 5331, 13916, 190, 177, 224), va(-1192, 11543, 9976, 127, 231, 199), va(-1192, 9115, 13218, 127, 220, 213), va(-1198, 6446, 15615, 127, 187, 238), va(-7838, 10585, 8500, 68, 223, 186), 
		va(-8548, 8054, 11579, 65, 211, 199), va(-8832, 5343, 13916, 63, 177, 224), va(-12513, 8042, 4584, 25, 199, 149), va(-13718, 5247, 7247, 20, 186, 161), va(-14200, 2421, 9422, 17, 152, 185), va(-14278, 4422, -988, 9, 167, 100), va(-15670, 1241, 1084, 3, 153, 109), va(-16230, -1735, 3018, 0, 118, 132), va(-12519, 795, -6560, 25, 135, 51), va(-13724, -2771, -5084, 20, 119, 58), 
		va(-14206, -5898, -3385, 17, 83, 79), va(-7850, -1753, -10476, 68, 112, 15), va(-8561, -5590, -9416, 65, 95, 20), va(-8844, -8826, -7886, 63, 58, 40), va(-1204, -2717, -11952, 126, 103, 2), va(-1204, -6657, -11049, 126, 86, 6), va(-1210, -9940, -9585, 126, 49, 26), va(5446, -1759, -10476, 185, 111, 15), va(6151, -5602, -9416, 188, 95, 20), va(6428, -8838, -7886, 190, 58, 40), 
		va(10115, 783, -6560, 228, 135, 51), va(11314, -2789, -5084, 233, 119, 58), va(11796, -5916, -3385, 236, 83, 79), va(10958, -240, 10549, 221, 102, 208), va(12850, -4138, 4566, 236, 72, 162), va(9392, -2283, 10784, 204, 75, 213), va(11037, -5675, 5566, 216, 51, 175), va(8548, -3355, 10892, 204, 75, 213), va(10067, -6482, 6090, 216, 51, 176), va(5940, 2494, 14760, 181, 124, 241), 
		va(5018, 102, 14447, 171, 94, 241), va(4524, -1162, 14266, 171, 93, 241), va(-1198, 3530, 16344, 127, 132, 253), va(-1198, 1006, 15832, 126, 100, 251), va(-1198, -331, 15537, 126, 100, 251), va(-8338, 2506, 14760, 72, 124, 241), va(-7422, 114, 14447, 82, 94, 241), va(-6928, -1150, 14266, 82, 93, 241), va(-13362, -228, 10549, 32, 102, 208), va(-11796, -2265, 10784, 49, 76, 213), 
		va(-10952, -3343, 10892, 49, 75, 213), va(-15260, -4114, 4566, 17, 72, 162), va(-13453, -5657, 5566, 37, 51, 175), va(-12477, -6464, 6090, 37, 51, 176), va(-13368, -8012, -1421, 32, 42, 116), va(-11802, -9049, 349, 49, 27, 138), va(-10958, -9585, 1289, 49, 27, 138), va(-8350, -10747, -5633, 72, 21, 83), va(-7434, -11434, -3319, 82, 9, 110), va(-6934, -11784, -2084, 82, 9, 111), 
		va(-1210, -11784, -7217, 126, 13, 70), va(-1210, -12338, -4699, 126, 2, 100), va(-1210, -12615, -3361, 126, 2, 101), va(5934, -10760, -5633, 181, 20, 83), va(5012, -11446, -3319, 171, 9, 110), va(4518, -11790, -2084, 171, 9, 111), va(10952, -8030, -1421, 221, 42, 116), va(9386, -9067, 349, 204, 27, 138), va(8542, -9603, 1289, 204, 26, 138), va(8079, -3964, 10952, 180, 50, 213), 
		va(9524, -6934, 6386, 188, 33, 187), va(5440, -5157, 9886, 136, 23, 200), va(6476, -7283, 6615, 138, 20, 195), va(-1204, -7416, 6705, 126, 20, 196), va(4247, -1873, 14163, 157, 62, 232), va(2699, -3656, 12181, 132, 26, 204), va(-1204, -1078, 15380, 126, 67, 239), va(-1204, -3090, 13049, 126, 27, 205), va(-6651, -1861, 14163, 96, 62, 232), va(-5108, -3650, 12181, 121, 26, 204), 
		va(-10488, -3946, 10952, 73, 50, 213), va(-7850, -5145, 9886, 117, 23, 200), va(-11934, -6922, 6386, 65, 33, 187), va(-8886, -7271, 6615, 115, 20, 195), va(-10488, -9892, 1813, 73, 17, 161), va(-7856, -9398, 3337, 117, 17, 191), va(-6663, -11983, -1397, 96, 4, 142), va(-5114, -10898, 1042, 121, 15, 187), va(-1210, -12772, -2608, 126, 0, 135), va(-1210, -11464, 174, 126, 14, 186), 
		va(4241, -11989, -1397, 157, 4, 142), va(2693, -10904, 1042, 132, 15, 187), va(8073, -9904, 1813, 180, 17, 161), va(5440, -9410, 3337, 136, 17, 191), va(-13218, 5349, -1590, 128, 20, 196), va(-13025, 6536, -566, 128, 133, 253), va(-17965, 6470, -524, 134, 122, 253), va(-17700, 5301, -1554, 137, 20, 195), va(-21019, 6012, -222, 159, 147, 247), va(-20513, 4934, -1319, 186, 32, 186), 
		va(-22068, 4759, 590, 181, 180, 228), va(-21483, 3940, -668, 250, 101, 141), va(-12663, 7217, -1012, 125, 251, 152), va(-18459, 7133, -951, 118, 246, 167), va(-21971, 6494, -536, 79, 237, 168), va(-23152, 4759, 590, 45, 189, 201), va(-12464, 6765, -2512, 124, 233, 57), va(-18730, 6663, -2446, 110, 232, 58), va(-22483, 5934, -1964, 47, 210, 73), va(-23743, 3940, -668, 0, 138, 120), 
		va(-12663, 5578, -3530, 125, 154, 2), va(-18465, 5494, -3476, 118, 138, 0), va(-21977, 4855, -3054, 79, 132, 9), va(-23158, 3120, -1927, 45, 82, 39), va(-13025, 4898, -3090, 127, 13, 69), va(-17965, 4831, -3048, 133, 9, 80), va(-21025, 4373, -2747, 160, 24, 60), va(-22068, 3120, -1927, 182, 57, 36), va(-21447, 2723, 1915, 186, 210, 202), va(-20959, 2150, 494, 242, 170, 97), 
		va(-19483, 506, 3355, 174, 226, 189), va(-19260, 48, 1855, 217, 200, 77), va(-16037, -1409, 4596, 155, 225, 201), va(-16230, -1735, 3018, 198, 213, 68), va(-22363, 2259, 2217, 57, 150, 230), va(-19899, -168, 3789, 75, 129, 242), va(-15676, -2319, 5187, 71, 88, 234), va(-22851, 1192, 1114, 15, 76, 160), va(-20128, -1349, 2765, 46, 45, 181), va(-15483, -3626, 4247, 62, 35, 186), 
		va(-22363, 620, -307, 57, 42, 62), va(-19905, -1807, 1271, 75, 22, 76), va(-15676, -3958, 2668, 73, 12, 117), va(-21447, 1084, -608, 187, 91, 20), va(-19489, -1132, 831, 175, 111, 10), va(-16037, -3048, 2078, 155, 99, 6), va(11573, 1548, 867, 86, 227, 60), va(11573, 2006, 4512, 116, 233, 194), va(16380, 3367, 2988, 108, 233, 193), va(15862, 2723, 102, 41, 205, 76), 
		va(17959, 5904, 162, 69, 224, 184), va(17308, 5259, -1542, 17, 182, 94), va(20260, 8368, -2078, 86, 238, 171), va(19092, 7687, -3126, 36, 204, 82), va(11573, -500, 6139, 174, 116, 244), va(17344, 1765, 4030, 196, 141, 232), va(19164, 5307, 548, 192, 170, 226), va(22429, 8368, -2078, 167, 177, 236), va(11567, -3644, 4247, 190, 34, 187), va(17863, -608, 2265, 222, 56, 172), 
		va(19815, 4012, -735, 238, 74, 158), va(23598, 7681, -3126, 199, 38, 181), va(11567, -4102, 596, 174, 15, 88), va(17338, -1253, -620, 197, 37, 70), va(19164, 3361, -2439, 192, 52, 47), va(22429, 7000, -4175, 167, 44, 39), va(11573, -1596, -1030, 119, 108, 1), va(16380, 343, -1662, 110, 109, 2), va(17959, 3958, -2831, 71, 110, 13), va(20260, 7006, -4175, 89, 129, 5), 
		va(21032, 8639, -2409, 114, 253, 133), va(19790, 8000, -3331, 82, 227, 64), va(21212, 8512, -2614, 133, 175, 9), va(20152, 8000, -3331, 209, 208, 75), va(20622, 8097, -2494, 188, 29, 73), va(19845, 7687, -3126, 223, 58, 173), va(23333, 8687, -2439, 189, 216, 191), va(23188, 8579, -2656, 110, 222, 44), va(22068, 8097, -2494, 113, 116, 1), va(24574, 8103, -3397, 252, 141, 115), 
		va(24255, 8127, -3415, 126, 232, 56), va(22851, 7687, -3126, 81, 226, 61), va(23333, 7464, -4319, 192, 103, 20), va(23188, 7615, -4132, 110, 241, 73), va(22068, 7277, -3753, 115, 236, 189), va(21025, 7416, -4289, 115, 172, 8), va(21212, 7554, -4090, 133, 253, 128), va(20622, 7277, -3753, 188, 128, 237), va(-1192, 12428, -6199, 127, 233, 57), va(1168, 12657, -4693, 231, 194, 154), 
		va(1536, 11898, -5855, 247, 161, 104), va(349, 11241, -4343, 227, 115, 203), va(590, 10747, -5102, 243, 84, 154), va(108, 10006, -3717, 217, 216, 130), va(307, 9591, -4355, 231, 187, 87), va(198, 13187, -3873, 187, 218, 191), va(-289, 11585, -3813, 184, 138, 239), va(-427, 10302, -3265, 179, 237, 163), va(-1192, 13386, -3566, 127, 227, 205), va(-1192, 11717, -3614, 127, 147, 252), 
		va(-1192, 10410, -3096, 127, 244, 174), va(-2578, 13187, -3873, 67, 218, 191), va(-2096, 11585, -3813, 69, 138, 239), va(-1958, 10302, -3265, 75, 237, 163), va(-3554, 12663, -4693, 22, 194, 154), va(-2735, 11241, -4343, 26, 115, 203), va(-2494, 10006, -3717, 36, 216, 130), va(-3922, 11904, -5855, 6, 161, 104), va(-2976, 10747, -5102, 10, 84, 154), va(-2699, 9591, -4355, 22, 187, 87), 
		va(-3554, 11145, -7018, 22, 128, 54), va(-2735, 10253, -5867, 26, 52, 106), va(-2494, 9175, -4994, 36, 159, 43), va(-2584, 10615, -7838, 66, 104, 17), va(-2102, 9910, -6398, 69, 29, 70), va(-1958, 8886, -5446, 75, 138, 11), va(-1192, 10416, -8145, 126, 96, 3), va(-1192, 9777, -6596, 126, 20, 57), va(-1192, 8771, -5614, 127, 130, 0), va(192, 10615, -7838, 186, 104, 17), 
		va(-289, 9904, -6398, 184, 29, 70), va(-433, 8880, -5446, 178, 138, 11), va(1168, 11145, -7018, 231, 128, 54), va(349, 10253, -5867, 227, 52, 106), va(108, 9175, -4994, 217, 159, 43), va(2536, 10085, -2060, 150, 238, 70), va(3120, 8886, -3897, 153, 231, 59), va(5693, 10603, -192, 161, 238, 77), va(6765, 8398, -3578, 166, 228, 61), va(7259, 10404, 1036, 173, 238, 86), 
		va(8573, 7693, -3126, 180, 223, 64), va(1000, 10922, -771, 140, 243, 78), va(2849, 12151, 2192, 146, 246, 89), va(3771, 12302, 3958, 153, 248, 102), va(-1192, 11241, -283, 127, 245, 81), va(-1192, 12742, 3090, 127, 249, 94), va(-1192, 13025, 5066, 127, 252, 108), va(-3385, 10928, -771, 113, 243, 78), va(-5235, 12157, 2192, 107, 246, 89), va(-6157, 12314, 3958, 100, 248, 102), 
		va(-4928, 10091, -2060, 103, 238, 70), va(-8079, 10609, -192, 92, 238, 77), va(-9645, 10416, 1036, 81, 238, 86), va(-5506, 8898, -3897, 100, 231, 59), va(-9151, 8410, -3578, 87, 228, 61), va(-10964, 7711, -3126, 73, 223, 64), va(-4928, 7699, -5735, 103, 223, 48), va(-8085, 6205, -6970, 92, 217, 44), va(-9651, 5000, -7289, 81, 209, 41), va(-3385, 6862, -7030, 113, 218, 39), 
		va(-5241, 4651, -9356, 107, 209, 32), va(-6163, 3102, -10211, 100, 198, 25), va(-1198, 6542, -7518, 127, 216, 36), va(-1198, 4066, -10253, 127, 206, 28), va(-1198, 2379, -11314, 127, 194, 19), va(994, 6856, -7030, 140, 218, 39), va(2849, 4644, -9356, 146, 209, 32), va(3765, 3090, -10211, 153, 198, 25), va(2536, 7693, -5735, 150, 223, 48), va(5687, 6193, -6970, 161, 217, 44), 
		va(7253, 4988, -7289, 173, 209, 41)
	);

	constant indices : indices_arr_t(0 to 575) := (
		idx(0, 1, 2), idx(2, 3, 0), 
		idx(3, 2, 4), idx(4, 5, 3), idx(5, 4, 6), idx(6, 7, 5), idx(1, 8, 9), idx(9, 2, 1), idx(2, 9, 10), idx(10, 4, 2), idx(4, 10, 11), idx(11, 6, 4), 
		idx(8, 12, 13), idx(13, 9, 8), idx(9, 13, 14), idx(14, 10, 9), idx(10, 14, 15), idx(15, 11, 10), idx(12, 16, 17), idx(17, 13, 12), idx(13, 17, 18), idx(18, 14, 13), 
		idx(14, 18, 19), idx(19, 15, 14), idx(16, 20, 21), idx(21, 17, 16), idx(17, 21, 22), idx(22, 18, 17), idx(18, 22, 23), idx(23, 19, 18), idx(20, 24, 25), idx(25, 21, 20), 
		idx(21, 25, 26), idx(26, 22, 21), idx(22, 26, 27), idx(27, 23, 22), idx(24, 28, 29), idx(29, 25, 24), idx(25, 29, 30), idx(30, 26, 25), idx(26, 30, 31), idx(31, 27, 26), 
		idx(28, 32, 33), idx(33, 29, 28), idx(29, 33, 34), idx(34, 30, 29), idx(30, 34, 35), idx(35, 31, 30), idx(32, 36, 37), idx(37, 33, 32), idx(33, 37, 38), idx(38, 34, 33), 
		idx(34, 38, 39), idx(39, 35, 34), idx(36, 40, 41), idx(41, 37, 36), idx(37, 41, 42), idx(42, 38, 37), idx(38, 42, 43), idx(43, 39, 38), idx(40, 44, 45), idx(45, 41, 40), 
		idx(41, 45, 46), idx(46, 42, 41), idx(42, 46, 47), idx(47, 43, 42), idx(44, 0, 3), idx(3, 45, 44), idx(45, 3, 5), idx(5, 46, 45), idx(46, 5, 7), idx(7, 47, 46), 
		idx(7, 6, 48), idx(48, 49, 7), idx(49, 48, 50), idx(50, 51, 49), idx(51, 50, 52), idx(52, 53, 51), idx(6, 11, 54), idx(54, 48, 6), idx(48, 54, 55), idx(55, 50, 48), 
		idx(50, 55, 56), idx(56, 52, 50), idx(11, 15, 57), idx(57, 54, 11), idx(54, 57, 58), idx(58, 55, 54), idx(55, 58, 59), idx(59, 56, 55), idx(15, 19, 60), idx(60, 57, 15), 
		idx(57, 60, 61), idx(61, 58, 57), idx(58, 61, 62), idx(62, 59, 58), idx(19, 23, 63), idx(63, 60, 19), idx(60, 63, 64), idx(64, 61, 60), idx(61, 64, 65), idx(65, 62, 61), 
		idx(23, 27, 66), idx(66, 63, 23), idx(63, 66, 67), idx(67, 64, 63), idx(64, 67, 68), idx(68, 65, 64), idx(27, 31, 69), idx(69, 66, 27), idx(66, 69, 70), idx(70, 67, 66), 
		idx(67, 70, 71), idx(71, 68, 67), idx(31, 35, 72), idx(72, 69, 31), idx(69, 72, 73), idx(73, 70, 69), idx(70, 73, 74), idx(74, 71, 70), idx(35, 39, 75), idx(75, 72, 35), 
		idx(72, 75, 76), idx(76, 73, 72), idx(73, 76, 77), idx(77, 74, 73), idx(39, 43, 78), idx(78, 75, 39), idx(75, 78, 79), idx(79, 76, 75), idx(76, 79, 80), idx(80, 77, 76), 
		idx(43, 47, 81), idx(81, 78, 43), idx(78, 81, 82), idx(82, 79, 78), idx(79, 82, 83), idx(83, 80, 79), idx(47, 7, 49), idx(49, 81, 47), idx(81, 49, 51), idx(51, 82, 81), 
		idx(82, 51, 53), idx(53, 83, 82), idx(53, 52, 84), idx(84, 85, 53), idx(85, 84, 86), idx(86, 87, 85), idx(87, 86, 88), idx(88, 89, 87), idx(52, 56, 90), idx(90, 84, 52), 
		idx(84, 90, 91), idx(91, 86, 84), idx(86, 91, 92), idx(92, 88, 86), idx(56, 59, 93), idx(93, 90, 56), idx(90, 93, 94), idx(94, 91, 90), idx(91, 94, 95), idx(95, 92, 91), 
		idx(59, 62, 96), idx(96, 93, 59), idx(93, 96, 97), idx(97, 94, 93), idx(94, 97, 98), idx(98, 95, 94), idx(62, 65, 99), idx(99, 96, 62), idx(96, 99, 100), idx(100, 97, 96), 
		idx(97, 100, 101), idx(101, 98, 97), idx(65, 68, 102), idx(102, 99, 65), idx(99, 102, 103), idx(103, 100, 99), idx(100, 103, 104), idx(104, 101, 100), idx(68, 71, 105), idx(105, 102, 68), 
		idx(102, 105, 106), idx(106, 103, 102), idx(103, 106, 107), idx(107, 104, 103), idx(71, 74, 108), idx(108, 105, 71), idx(105, 108, 109), idx(109, 106, 105), idx(106, 109, 110), idx(110, 107, 106), 
		idx(74, 77, 111), idx(111, 108, 74), idx(108, 111, 112), idx(112, 109, 108), idx(109, 112, 113), idx(113, 110, 109), idx(77, 80, 114), idx(114, 111, 77), idx(111, 114, 115), idx(115, 112, 111), 
		idx(112, 115, 116), idx(116, 113, 112), idx(80, 83, 117), idx(117, 114, 80), idx(114, 117, 118), idx(118, 115, 114), idx(115, 118, 119), idx(119, 116, 115), idx(83, 53, 85), idx(85, 117, 83), 
		idx(117, 85, 87), idx(87, 118, 117), idx(118, 87, 89), idx(89, 119, 118), idx(89, 88, 120), idx(120, 121, 89), idx(121, 120, 122), idx(122, 123, 121), idx(123, 122, 124), idx(124, 124, 123), 
		idx(88, 92, 125), idx(125, 120, 88), idx(120, 125, 126), idx(126, 122, 120), idx(122, 126, 124), idx(124, 124, 122), idx(92, 95, 127), idx(127, 125, 92), idx(125, 127, 128), idx(128, 126, 125), 
		idx(126, 128, 124), idx(124, 124, 126), idx(95, 98, 129), idx(129, 127, 95), idx(127, 129, 130), idx(130, 128, 127), idx(128, 130, 124), idx(124, 124, 128), idx(98, 101, 131), idx(131, 129, 98), 
		idx(129, 131, 132), idx(132, 130, 129), idx(130, 132, 124), idx(124, 124, 130), idx(101, 104, 133), idx(133, 131, 101), idx(131, 133, 134), idx(134, 132, 131), idx(132, 134, 124), idx(124, 124, 132), 
		idx(104, 107, 135), idx(135, 133, 104), idx(133, 135, 136), idx(136, 134, 133), idx(134, 136, 124), idx(124, 124, 134), idx(107, 110, 137), idx(137, 135, 107), idx(135, 137, 138), idx(138, 136, 135), 
		idx(136, 138, 124), idx(124, 124, 136), idx(110, 113, 139), idx(139, 137, 110), idx(137, 139, 140), idx(140, 138, 137), idx(138, 140, 124), idx(124, 124, 138), idx(113, 116, 141), idx(141, 139, 113), 
		idx(139, 141, 142), idx(142, 140, 139), idx(140, 142, 124), idx(124, 124, 140), idx(116, 119, 143), idx(143, 141, 116), idx(141, 143, 144), idx(144, 142, 141), idx(142, 144, 124), idx(124, 124, 142), 
		idx(119, 89, 121), idx(121, 143, 119), idx(143, 121, 123), idx(123, 144, 143), idx(144, 123, 124), idx(124, 124, 144), idx(145, 146, 147), idx(147, 148, 145), idx(148, 147, 149), idx(149, 150, 148), 
		idx(150, 149, 151), idx(151, 152, 150), idx(146, 153, 154), idx(154, 147, 146), idx(147, 154, 155), idx(155, 149, 147), idx(149, 155, 156), idx(156, 151, 149), idx(153, 157, 158), idx(158, 154, 153), 
		idx(154, 158, 159), idx(159, 155, 154), idx(155, 159, 160), idx(160, 156, 155), idx(157, 161, 162), idx(162, 158, 157), idx(158, 162, 163), idx(163, 159, 158), idx(159, 163, 164), idx(164, 160, 159), 
		idx(161, 165, 166), idx(166, 162, 161), idx(162, 166, 167), idx(167, 163, 162), idx(163, 167, 168), idx(168, 164, 163), idx(165, 145, 148), idx(148, 166, 165), idx(166, 148, 150), idx(150, 167, 166), 
		idx(167, 150, 152), idx(152, 168, 167), idx(152, 151, 169), idx(169, 170, 152), idx(170, 169, 171), idx(171, 172, 170), idx(172, 171, 173), idx(173, 174, 172), idx(151, 156, 175), idx(175, 169, 151), 
		idx(169, 175, 176), idx(176, 171, 169), idx(171, 176, 177), idx(177, 173, 171), idx(156, 160, 178), idx(178, 175, 156), idx(175, 178, 179), idx(179, 176, 175), idx(176, 179, 180), idx(180, 177, 176), 
		idx(160, 164, 181), idx(181, 178, 160), idx(178, 181, 182), idx(182, 179, 178), idx(179, 182, 183), idx(183, 180, 179), idx(164, 168, 184), idx(184, 181, 164), idx(181, 184, 185), idx(185, 182, 181), 
		idx(182, 185, 186), idx(186, 183, 182), idx(168, 152, 170), idx(170, 184, 168), idx(184, 170, 172), idx(172, 185, 184), idx(185, 172, 174), idx(174, 186, 185), idx(187, 188, 189), idx(189, 190, 187), 
		idx(190, 189, 191), idx(191, 192, 190), idx(192, 191, 193), idx(193, 194, 192), idx(188, 195, 196), idx(196, 189, 188), idx(189, 196, 197), idx(197, 191, 189), idx(191, 197, 198), idx(198, 193, 191), 
		idx(195, 199, 200), idx(200, 196, 195), idx(196, 200, 201), idx(201, 197, 196), idx(197, 201, 202), idx(202, 198, 197), idx(199, 203, 204), idx(204, 200, 199), idx(200, 204, 205), idx(205, 201, 200), 
		idx(201, 205, 206), idx(206, 202, 201), idx(203, 207, 208), idx(208, 204, 203), idx(204, 208, 209), idx(209, 205, 204), idx(205, 209, 210), idx(210, 206, 205), idx(207, 187, 190), idx(190, 208, 207), 
		idx(208, 190, 192), idx(192, 209, 208), idx(209, 192, 194), idx(194, 210, 209), idx(194, 193, 211), idx(211, 212, 194), idx(212, 211, 213), idx(213, 214, 212), idx(214, 213, 215), idx(215, 216, 214), 
		idx(193, 198, 217), idx(217, 211, 193), idx(211, 217, 218), idx(218, 213, 211), idx(213, 218, 219), idx(219, 215, 213), idx(198, 202, 220), idx(220, 217, 198), idx(217, 220, 221), idx(221, 218, 217), 
		idx(218, 221, 222), idx(222, 219, 218), idx(202, 206, 223), idx(223, 220, 202), idx(220, 223, 224), idx(224, 221, 220), idx(221, 224, 225), idx(225, 222, 221), idx(206, 210, 226), idx(226, 223, 206), 
		idx(223, 226, 227), idx(227, 224, 223), idx(224, 227, 228), idx(228, 225, 224), idx(210, 194, 212), idx(212, 226, 210), idx(226, 212, 214), idx(214, 227, 226), idx(227, 214, 216), idx(216, 228, 227), 
		idx(229, 229, 230), idx(230, 231, 229), idx(231, 230, 232), idx(232, 233, 231), idx(233, 232, 234), idx(234, 235, 233), idx(229, 229, 236), idx(236, 230, 229), idx(230, 236, 237), idx(237, 232, 230), 
		idx(232, 237, 238), idx(238, 234, 232), idx(229, 229, 239), idx(239, 236, 229), idx(236, 239, 240), idx(240, 237, 236), idx(237, 240, 241), idx(241, 238, 237), idx(229, 229, 242), idx(242, 239, 229), 
		idx(239, 242, 243), idx(243, 240, 239), idx(240, 243, 244), idx(244, 241, 240), idx(229, 229, 245), idx(245, 242, 229), idx(242, 245, 246), idx(246, 243, 242), idx(243, 246, 247), idx(247, 244, 243), 
		idx(229, 229, 248), idx(248, 245, 229), idx(245, 248, 249), idx(249, 246, 245), idx(246, 249, 250), idx(250, 247, 246), idx(229, 229, 251), idx(251, 248, 229), idx(248, 251, 252), idx(252, 249, 248), 
		idx(249, 252, 253), idx(253, 250, 249), idx(229, 229, 254), idx(254, 251, 229), idx(251, 254, 255), idx(255, 252, 251), idx(252, 255, 256), idx(256, 253, 252), idx(229, 229, 257), idx(257, 254, 229), 
		idx(254, 257, 258), idx(258, 255, 254), idx(255, 258, 259), idx(259, 256, 255), idx(229, 229, 260), idx(260, 257, 229), idx(257, 260, 261), idx(261, 258, 257), idx(258, 261, 262), idx(262, 259, 258), 
		idx(229, 229, 263), idx(263, 260, 229), idx(260, 263, 264), idx(264, 261, 260), idx(261, 264, 265), idx(265, 262, 261), idx(229, 229, 231), idx(231, 263, 229), idx(263, 231, 233), idx(233, 264, 263), 
		idx(264, 233, 235), idx(235, 265, 264), idx(235, 234, 266), idx(266, 267, 235), idx(267, 266, 268), idx(268, 269, 267), idx(269, 268, 270), idx(270, 271, 269), idx(234, 238, 272), idx(272, 266, 234), 
		idx(266, 272, 273), idx(273, 268, 266), idx(268, 273, 274), idx(274, 270, 268), idx(238, 241, 275), idx(275, 272, 238), idx(272, 275, 276), idx(276, 273, 272), idx(273, 276, 277), idx(277, 274, 273), 
		idx(241, 244, 278), idx(278, 275, 241), idx(275, 278, 279), idx(279, 276, 275), idx(276, 279, 280), idx(280, 277, 276), idx(244, 247, 281), idx(281, 278, 244), idx(278, 281, 282), idx(282, 279, 278), 
		idx(279, 282, 283), idx(283, 280, 279), idx(247, 250, 284), idx(284, 281, 247), idx(281, 284, 285), idx(285, 282, 281), idx(282, 285, 286), idx(286, 283, 282), idx(250, 253, 287), idx(287, 284, 250), 
		idx(284, 287, 288), idx(288, 285, 284), idx(285, 288, 289), idx(289, 286, 285), idx(253, 256, 290), idx(290, 287, 253), idx(287, 290, 291), idx(291, 288, 287), idx(288, 291, 292), idx(292, 289, 288), 
		idx(256, 259, 293), idx(293, 290, 256), idx(290, 293, 294), idx(294, 291, 290), idx(291, 294, 295), idx(295, 292, 291), idx(259, 262, 296), idx(296, 293, 259), idx(293, 296, 297), idx(297, 294, 293), 
		idx(294, 297, 298), idx(298, 295, 294), idx(262, 265, 299), idx(299, 296, 262), idx(296, 299, 300), idx(300, 297, 296), idx(297, 300, 301), idx(301, 298, 297), idx(265, 235, 267), idx(267, 299, 265), 
		idx(299, 267, 269), idx(269, 300, 299), idx(300, 269, 271), idx(271, 301, 300)
	);

end package renderer_mesh;
