use work.common.all;

package renderer_mesh is
	constant vertices : vertex_arr_3d_t(0 to 528) := (
		point3d(206, 135, 79), point3d(216, 102, 79), point3d(218, 102, 72), point3d(207, 135, 72), point3d(216, 102, 69), point3d(205, 135, 69), point3d(212, 101, 72), point3d(201, 135, 72), point3d(207, 100, 79), point3d(196, 135, 79), point3d(245, 75, 79), 
		point3d(246, 76, 72), point3d(244, 75, 69), point3d(241, 73, 72), point3d(238, 71, 79), point3d(288, 58, 79), point3d(288, 59, 72), point3d(287, 57, 69), point3d(286, 55, 72), point3d(284, 52, 79), point3d(340, 51, 79), 
		point3d(340, 52, 72), point3d(340, 51, 69), point3d(340, 48, 72), point3d(340, 45, 79), point3d(397, 58, 79), point3d(394, 59, 72), point3d(394, 57, 69), point3d(395, 55, 72), point3d(397, 52, 79), point3d(439, 75, 79), 
		point3d(436, 76, 72), point3d(437, 75, 69), point3d(440, 73, 72), point3d(443, 71, 79), point3d(466, 102, 79), point3d(464, 102, 72), point3d(465, 102, 69), point3d(469, 101, 72), point3d(474, 100, 79), point3d(475, 135, 79), 
		point3d(473, 135, 72), point3d(476, 135, 69), point3d(480, 135, 72), point3d(485, 135, 79), point3d(465, 168, 79), point3d(463, 167, 72), point3d(465, 168, 69), point3d(469, 169, 72), point3d(474, 170, 79), point3d(436, 194, 79), 
		point3d(435, 193, 72), point3d(436, 194, 69), point3d(440, 196, 72), point3d(443, 199, 79), point3d(393, 212, 79), point3d(393, 211, 72), point3d(394, 212, 69), point3d(395, 215, 72), point3d(397, 218, 79), point3d(340, 219, 79), 
		point3d(340, 217, 72), point3d(340, 219, 69), point3d(340, 222, 72), point3d(340, 225, 79), point3d(288, 212, 79), point3d(288, 211, 72), point3d(287, 212, 69), point3d(286, 215, 72), point3d(284, 218, 79), point3d(245, 194, 79), 
		point3d(246, 193, 72), point3d(244, 194, 69), point3d(241, 196, 72), point3d(238, 199, 79), point3d(216, 168, 79), point3d(218, 167, 72), point3d(216, 168, 69), point3d(212, 169, 72), point3d(207, 170, 79), point3d(191, 95, 115), 
		point3d(178, 135, 115), point3d(177, 92, 150), point3d(163, 135, 150), point3d(167, 89, 184), point3d(152, 135, 184), point3d(163, 88, 217), point3d(148, 135, 217), point3d(225, 63, 115), point3d(214, 56, 150), point3d(207, 52, 184), 
		point3d(204, 50, 217), point3d(277, 42, 115), point3d(271, 33, 150), point3d(266, 27, 184), point3d(265, 24, 217), point3d(340, 34, 115), point3d(340, 24, 150), point3d(340, 18, 184), point3d(340, 15, 217), point3d(404, 42, 115), 
		point3d(410, 33, 150), point3d(414, 27, 184), point3d(416, 24, 217), point3d(456, 63, 115), point3d(467, 56, 150), point3d(474, 52, 184), point3d(477, 50, 217), point3d(490, 95, 115), point3d(504, 92, 150), point3d(514, 89, 184), 
		point3d(518, 88, 217), point3d(503, 135, 115), point3d(518, 135, 150), point3d(529, 135, 184), point3d(533, 135, 217), point3d(490, 174, 115), point3d(504, 178, 150), point3d(514, 181, 184), point3d(518, 182, 217), point3d(456, 206, 115), 
		point3d(467, 213, 150), point3d(474, 218, 184), point3d(477, 220, 217), point3d(404, 228, 115), point3d(410, 237, 150), point3d(414, 243, 184), point3d(416, 245, 217), point3d(340, 236, 115), point3d(340, 245, 150), point3d(340, 252, 184), 
		point3d(340, 255, 217), point3d(277, 228, 115), point3d(271, 237, 150), point3d(266, 243, 184), point3d(265, 245, 217), point3d(225, 206, 115), point3d(214, 213, 150), point3d(207, 218, 184), point3d(204, 220, 217), point3d(191, 174, 115), 
		point3d(177, 178, 150), point3d(167, 181, 184), point3d(163, 182, 217), point3d(170, 90, 244), point3d(155, 135, 244), point3d(185, 94, 264), point3d(172, 135, 264), point3d(200, 98, 278), point3d(188, 135, 278), point3d(207, 100, 286), 
		point3d(196, 135, 286), point3d(209, 53, 244), point3d(221, 60, 264), point3d(233, 68, 278), point3d(238, 71, 286), point3d(268, 29, 244), point3d(274, 38, 264), point3d(281, 48, 278), point3d(284, 52, 286), point3d(340, 20, 244), 
		point3d(340, 30, 264), point3d(340, 40, 278), point3d(340, 45, 286), point3d(413, 29, 244), point3d(407, 38, 264), point3d(400, 48, 278), point3d(397, 52, 286), point3d(472, 53, 244), point3d(460, 60, 264), point3d(448, 68, 278), 
		point3d(443, 71, 286), point3d(511, 90, 244), point3d(496, 94, 264), point3d(481, 98, 278), point3d(474, 100, 286), point3d(526, 135, 244), point3d(509, 135, 264), point3d(493, 135, 278), point3d(485, 135, 286), point3d(511, 180, 244), 
		point3d(496, 176, 264), point3d(481, 172, 278), point3d(474, 170, 286), point3d(472, 216, 244), point3d(460, 209, 264), point3d(448, 202, 278), point3d(443, 199, 286), point3d(413, 241, 244), point3d(407, 231, 264), point3d(400, 222, 278), 
		point3d(397, 218, 286), point3d(340, 250, 244), point3d(340, 240, 264), point3d(340, 229, 278), point3d(340, 225, 286), point3d(268, 241, 244), point3d(274, 231, 264), point3d(281, 222, 278), point3d(284, 218, 286), point3d(209, 216, 244), 
		point3d(221, 209, 264), point3d(233, 202, 278), point3d(238, 199, 286), point3d(170, 180, 244), point3d(185, 176, 264), point3d(200, 172, 278), point3d(207, 170, 286), point3d(210, 100, 291), point3d(199, 135, 291), point3d(226, 105, 295), 
		point3d(217, 135, 295), point3d(266, 115, 298), point3d(260, 135, 298), point3d(340, 135, 300), point3d(240, 73, 291), point3d(253, 80, 295), point3d(283, 99, 298), point3d(285, 54, 291), point3d(292, 64, 295), point3d(309, 89, 298), 
		point3d(340, 47, 291), point3d(340, 58, 295), point3d(340, 85, 298), point3d(396, 54, 291), point3d(389, 64, 295), point3d(372, 89, 298), point3d(441, 73, 291), point3d(428, 80, 295), point3d(398, 99, 298), point3d(471, 100, 291), 
		point3d(455, 105, 295), point3d(415, 115, 298), point3d(482, 135, 291), point3d(464, 135, 295), point3d(421, 135, 298), point3d(471, 169, 291), point3d(455, 165, 295), point3d(415, 154, 298), point3d(441, 197, 291), point3d(428, 189, 295), 
		point3d(398, 170, 298), point3d(396, 216, 291), point3d(389, 206, 295), point3d(372, 181, 298), point3d(340, 223, 291), point3d(340, 212, 295), point3d(340, 185, 298), point3d(285, 216, 291), point3d(292, 206, 295), point3d(309, 181, 298), 
		point3d(240, 197, 291), point3d(253, 189, 295), point3d(283, 170, 298), point3d(210, 169, 291), point3d(226, 165, 295), point3d(266, 154, 298), point3d(495, 135, 113), point3d(493, 125, 110), point3d(541, 125, 110), point3d(540, 135, 113), 
		point3d(576, 125, 113), point3d(573, 135, 116), point3d(598, 125, 120), point3d(594, 135, 122), point3d(605, 125, 134), point3d(601, 135, 134), point3d(490, 121, 103), point3d(544, 121, 103), point3d(583, 121, 107), point3d(607, 121, 116), 
		point3d(615, 121, 134), point3d(486, 125, 96), point3d(547, 125, 96), point3d(590, 125, 100), point3d(616, 125, 112), point3d(625, 125, 134), point3d(485, 135, 92), point3d(548, 135, 93), point3d(593, 135, 98), point3d(620, 135, 110), 
		point3d(630, 135, 134), point3d(486, 145, 96), point3d(547, 145, 96), point3d(590, 145, 100), point3d(616, 145, 112), point3d(625, 145, 134), point3d(490, 148, 103), point3d(544, 148, 103), point3d(583, 148, 107), point3d(607, 148, 116), 
		point3d(615, 148, 134), point3d(493, 145, 110), point3d(541, 145, 110), point3d(576, 145, 113), point3d(598, 145, 120), point3d(605, 145, 134), point3d(601, 125, 154), point3d(597, 135, 153), point3d(588, 125, 178), point3d(585, 135, 175), 
		point3d(565, 125, 201), point3d(564, 135, 198), point3d(532, 125, 221), point3d(610, 121, 158), point3d(594, 121, 184), point3d(567, 121, 209), point3d(528, 121, 230), point3d(619, 125, 162), point3d(601, 125, 190), point3d(570, 125, 216), 
		point3d(525, 125, 240), point3d(623, 135, 164), point3d(604, 135, 193), point3d(571, 135, 220), point3d(524, 135, 244), point3d(619, 145, 162), point3d(601, 145, 190), point3d(570, 145, 216), point3d(525, 145, 240), point3d(610, 148, 158), 
		point3d(594, 148, 184), point3d(567, 148, 209), point3d(528, 148, 230), point3d(601, 145, 154), point3d(588, 145, 178), point3d(565, 145, 201), point3d(532, 145, 221), point3d(177, 135, 168), point3d(177, 113, 180), point3d(127, 115, 167), 
		point3d(130, 135, 158), point3d(106, 119, 139), point3d(110, 135, 134), point3d(94, 124, 106), point3d(99, 135, 104), point3d(71, 126, 79), point3d(80, 135, 79), point3d(177, 105, 206), point3d(119, 108, 186), point3d(96, 114, 150), 
		point3d(82, 121, 110), point3d(51, 124, 79), point3d(177, 113, 232), point3d(111, 115, 206), point3d(86, 119, 161), point3d(70, 124, 114), point3d(32, 126, 79), point3d(177, 135, 244), point3d(108, 135, 214), point3d(82, 135, 167), 
		point3d(64, 135, 116), point3d(23, 135, 79), point3d(177, 157, 232), point3d(111, 155, 206), point3d(86, 150, 161), point3d(70, 145, 114), point3d(32, 143, 79), point3d(177, 164, 206), point3d(119, 162, 186), point3d(96, 155, 150), 
		point3d(82, 149, 110), point3d(51, 146, 79), point3d(177, 157, 180), point3d(127, 155, 167), point3d(106, 150, 139), point3d(94, 145, 106), point3d(71, 143, 79), point3d(64, 127, 74), point3d(73, 135, 75), point3d(59, 128, 73), 
		point3d(68, 135, 73), point3d(59, 129, 74), point3d(67, 135, 75), point3d(65, 130, 79), point3d(71, 135, 79), point3d(42, 124, 74), point3d(39, 126, 72), point3d(42, 127, 74), point3d(51, 128, 79), point3d(21, 127, 74), 
		point3d(19, 128, 72), point3d(25, 129, 73), point3d(38, 130, 79), point3d(11, 135, 73), point3d(10, 135, 71), point3d(17, 135, 73), point3d(32, 135, 79), point3d(21, 143, 74), point3d(19, 142, 72), point3d(25, 140, 73), 
		point3d(38, 140, 79), point3d(42, 145, 74), point3d(39, 144, 72), point3d(42, 142, 74), point3d(51, 142, 79), point3d(64, 143, 74), point3d(59, 142, 73), point3d(59, 140, 74), point3d(65, 140, 79), point3d(340, 135, 9), 
		point3d(310, 127, 14), point3d(308, 135, 14), point3d(312, 127, 25), point3d(309, 135, 25), point3d(323, 130, 39), point3d(321, 135, 39), point3d(323, 130, 51), point3d(321, 135, 51), point3d(317, 120, 14), point3d(318, 121, 25), 
		point3d(327, 126, 39), point3d(327, 126, 51), point3d(328, 116, 14), point3d(328, 117, 25), point3d(333, 124, 39), point3d(333, 124, 51), point3d(340, 114, 14), point3d(340, 115, 25), point3d(340, 123, 39), point3d(340, 123, 51), 
		point3d(353, 116, 14), point3d(353, 117, 25), point3d(348, 124, 39), point3d(348, 124, 51), point3d(364, 120, 14), point3d(363, 121, 25), point3d(354, 126, 39), point3d(354, 126, 51), point3d(371, 127, 14), point3d(369, 127, 25), 
		point3d(358, 130, 39), point3d(358, 130, 51), point3d(373, 135, 14), point3d(372, 135, 25), point3d(359, 135, 39), point3d(360, 135, 51), point3d(371, 143, 14), point3d(369, 142, 25), point3d(358, 139, 39), point3d(358, 140, 51), 
		point3d(364, 149, 14), point3d(363, 149, 25), point3d(354, 143, 39), point3d(354, 143, 51), point3d(353, 154, 14), point3d(353, 153, 25), point3d(348, 146, 39), point3d(348, 146, 51), point3d(340, 155, 14), point3d(340, 154, 25), 
		point3d(340, 147, 39), point3d(340, 147, 51), point3d(328, 154, 14), point3d(328, 153, 25), point3d(333, 146, 39), point3d(333, 146, 51), point3d(317, 149, 14), point3d(318, 149, 25), point3d(327, 143, 39), point3d(327, 143, 51), 
		point3d(310, 143, 14), point3d(312, 142, 25), point3d(323, 139, 39), point3d(323, 140, 51), point3d(300, 124, 59), point3d(296, 135, 59), point3d(267, 115, 65), point3d(261, 135, 65), point3d(238, 108, 70), point3d(229, 135, 70), 
		point3d(225, 104, 79), point3d(215, 135, 79), point3d(309, 115, 59), point3d(284, 100, 65), point3d(261, 86, 70), point3d(252, 80, 79), point3d(323, 110, 59), point3d(309, 89, 65), point3d(297, 71, 70), point3d(291, 63, 79), 
		point3d(340, 108, 59), point3d(340, 85, 65), point3d(340, 66, 70), point3d(340, 57, 79), point3d(358, 110, 59), point3d(372, 89, 65), point3d(384, 71, 70), point3d(390, 63, 79), point3d(372, 115, 59), point3d(397, 100, 65), 
		point3d(420, 86, 70), point3d(429, 80, 79), point3d(381, 124, 59), point3d(414, 115, 65), point3d(443, 108, 70), point3d(456, 104, 79), point3d(384, 135, 59), point3d(420, 135, 65), point3d(452, 135, 70), point3d(466, 135, 79), 
		point3d(381, 146, 59), point3d(414, 154, 65), point3d(443, 162, 70), point3d(456, 165, 79), point3d(372, 154, 59), point3d(397, 170, 65), point3d(420, 184, 70), point3d(429, 190, 79), point3d(358, 160, 59), point3d(372, 180, 65), 
		point3d(384, 199, 70), point3d(390, 207, 79), point3d(340, 162, 59), point3d(340, 184, 65), point3d(340, 204, 70), point3d(340, 213, 79), point3d(323, 160, 59), point3d(309, 180, 65), point3d(297, 199, 70), point3d(291, 207, 79), 
		point3d(309, 154, 59), point3d(284, 170, 65), point3d(261, 184, 70), point3d(252, 190, 79), point3d(300, 146, 59), point3d(267, 154, 65), point3d(238, 162, 70), point3d(225, 165, 79)
	);

	constant indices : indices_arr_t(0 to 1023) := (
		idx(0, 1, 2), idx(2, 3, 0), 
		idx(3, 2, 4), idx(4, 5, 3), idx(5, 4, 6), idx(6, 7, 5), idx(7, 6, 8), idx(8, 9, 7), idx(1, 10, 11), idx(11, 2, 1), idx(2, 11, 12), idx(12, 4, 2), 
		idx(4, 12, 13), idx(13, 6, 4), idx(6, 13, 14), idx(14, 8, 6), idx(10, 15, 16), idx(16, 11, 10), idx(11, 16, 17), idx(17, 12, 11), idx(12, 17, 18), idx(18, 13, 12), 
		idx(13, 18, 19), idx(19, 14, 13), idx(15, 20, 21), idx(21, 16, 15), idx(16, 21, 22), idx(22, 17, 16), idx(17, 22, 23), idx(23, 18, 17), idx(18, 23, 24), idx(24, 19, 18), 
		idx(20, 25, 26), idx(26, 21, 20), idx(21, 26, 27), idx(27, 22, 21), idx(22, 27, 28), idx(28, 23, 22), idx(23, 28, 29), idx(29, 24, 23), idx(25, 30, 31), idx(31, 26, 25), 
		idx(26, 31, 32), idx(32, 27, 26), idx(27, 32, 33), idx(33, 28, 27), idx(28, 33, 34), idx(34, 29, 28), idx(30, 35, 36), idx(36, 31, 30), idx(31, 36, 37), idx(37, 32, 31), 
		idx(32, 37, 38), idx(38, 33, 32), idx(33, 38, 39), idx(39, 34, 33), idx(35, 40, 41), idx(41, 36, 35), idx(36, 41, 42), idx(42, 37, 36), idx(37, 42, 43), idx(43, 38, 37), 
		idx(38, 43, 44), idx(44, 39, 38), idx(40, 45, 46), idx(46, 41, 40), idx(41, 46, 47), idx(47, 42, 41), idx(42, 47, 48), idx(48, 43, 42), idx(43, 48, 49), idx(49, 44, 43), 
		idx(45, 50, 51), idx(51, 46, 45), idx(46, 51, 52), idx(52, 47, 46), idx(47, 52, 53), idx(53, 48, 47), idx(48, 53, 54), idx(54, 49, 48), idx(50, 55, 56), idx(56, 51, 50), 
		idx(51, 56, 57), idx(57, 52, 51), idx(52, 57, 58), idx(58, 53, 52), idx(53, 58, 59), idx(59, 54, 53), idx(55, 60, 61), idx(61, 56, 55), idx(56, 61, 62), idx(62, 57, 56), 
		idx(57, 62, 63), idx(63, 58, 57), idx(58, 63, 64), idx(64, 59, 58), idx(60, 65, 66), idx(66, 61, 60), idx(61, 66, 67), idx(67, 62, 61), idx(62, 67, 68), idx(68, 63, 62), 
		idx(63, 68, 69), idx(69, 64, 63), idx(65, 70, 71), idx(71, 66, 65), idx(66, 71, 72), idx(72, 67, 66), idx(67, 72, 73), idx(73, 68, 67), idx(68, 73, 74), idx(74, 69, 68), 
		idx(70, 75, 76), idx(76, 71, 70), idx(71, 76, 77), idx(77, 72, 71), idx(72, 77, 78), idx(78, 73, 72), idx(73, 78, 79), idx(79, 74, 73), idx(75, 0, 3), idx(3, 76, 75), 
		idx(76, 3, 5), idx(5, 77, 76), idx(77, 5, 7), idx(7, 78, 77), idx(78, 7, 9), idx(9, 79, 78), idx(9, 8, 80), idx(80, 81, 9), idx(81, 80, 82), idx(82, 83, 81), 
		idx(83, 82, 84), idx(84, 85, 83), idx(85, 84, 86), idx(86, 87, 85), idx(8, 14, 88), idx(88, 80, 8), idx(80, 88, 89), idx(89, 82, 80), idx(82, 89, 90), idx(90, 84, 82), 
		idx(84, 90, 91), idx(91, 86, 84), idx(14, 19, 92), idx(92, 88, 14), idx(88, 92, 93), idx(93, 89, 88), idx(89, 93, 94), idx(94, 90, 89), idx(90, 94, 95), idx(95, 91, 90), 
		idx(19, 24, 96), idx(96, 92, 19), idx(92, 96, 97), idx(97, 93, 92), idx(93, 97, 98), idx(98, 94, 93), idx(94, 98, 99), idx(99, 95, 94), idx(24, 29, 100), idx(100, 96, 24), 
		idx(96, 100, 101), idx(101, 97, 96), idx(97, 101, 102), idx(102, 98, 97), idx(98, 102, 103), idx(103, 99, 98), idx(29, 34, 104), idx(104, 100, 29), idx(100, 104, 105), idx(105, 101, 100), 
		idx(101, 105, 106), idx(106, 102, 101), idx(102, 106, 107), idx(107, 103, 102), idx(34, 39, 108), idx(108, 104, 34), idx(104, 108, 109), idx(109, 105, 104), idx(105, 109, 110), idx(110, 106, 105), 
		idx(106, 110, 111), idx(111, 107, 106), idx(39, 44, 112), idx(112, 108, 39), idx(108, 112, 113), idx(113, 109, 108), idx(109, 113, 114), idx(114, 110, 109), idx(110, 114, 115), idx(115, 111, 110), 
		idx(44, 49, 116), idx(116, 112, 44), idx(112, 116, 117), idx(117, 113, 112), idx(113, 117, 118), idx(118, 114, 113), idx(114, 118, 119), idx(119, 115, 114), idx(49, 54, 120), idx(120, 116, 49), 
		idx(116, 120, 121), idx(121, 117, 116), idx(117, 121, 122), idx(122, 118, 117), idx(118, 122, 123), idx(123, 119, 118), idx(54, 59, 124), idx(124, 120, 54), idx(120, 124, 125), idx(125, 121, 120), 
		idx(121, 125, 126), idx(126, 122, 121), idx(122, 126, 127), idx(127, 123, 122), idx(59, 64, 128), idx(128, 124, 59), idx(124, 128, 129), idx(129, 125, 124), idx(125, 129, 130), idx(130, 126, 125), 
		idx(126, 130, 131), idx(131, 127, 126), idx(64, 69, 132), idx(132, 128, 64), idx(128, 132, 133), idx(133, 129, 128), idx(129, 133, 134), idx(134, 130, 129), idx(130, 134, 135), idx(135, 131, 130), 
		idx(69, 74, 136), idx(136, 132, 69), idx(132, 136, 137), idx(137, 133, 132), idx(133, 137, 138), idx(138, 134, 133), idx(134, 138, 139), idx(139, 135, 134), idx(74, 79, 140), idx(140, 136, 74), 
		idx(136, 140, 141), idx(141, 137, 136), idx(137, 141, 142), idx(142, 138, 137), idx(138, 142, 143), idx(143, 139, 138), idx(79, 9, 81), idx(81, 140, 79), idx(140, 81, 83), idx(83, 141, 140), 
		idx(141, 83, 85), idx(85, 142, 141), idx(142, 85, 87), idx(87, 143, 142), idx(87, 86, 144), idx(144, 145, 87), idx(145, 144, 146), idx(146, 147, 145), idx(147, 146, 148), idx(148, 149, 147), 
		idx(149, 148, 150), idx(150, 151, 149), idx(86, 91, 152), idx(152, 144, 86), idx(144, 152, 153), idx(153, 146, 144), idx(146, 153, 154), idx(154, 148, 146), idx(148, 154, 155), idx(155, 150, 148), 
		idx(91, 95, 156), idx(156, 152, 91), idx(152, 156, 157), idx(157, 153, 152), idx(153, 157, 158), idx(158, 154, 153), idx(154, 158, 159), idx(159, 155, 154), idx(95, 99, 160), idx(160, 156, 95), 
		idx(156, 160, 161), idx(161, 157, 156), idx(157, 161, 162), idx(162, 158, 157), idx(158, 162, 163), idx(163, 159, 158), idx(99, 103, 164), idx(164, 160, 99), idx(160, 164, 165), idx(165, 161, 160), 
		idx(161, 165, 166), idx(166, 162, 161), idx(162, 166, 167), idx(167, 163, 162), idx(103, 107, 168), idx(168, 164, 103), idx(164, 168, 169), idx(169, 165, 164), idx(165, 169, 170), idx(170, 166, 165), 
		idx(166, 170, 171), idx(171, 167, 166), idx(107, 111, 172), idx(172, 168, 107), idx(168, 172, 173), idx(173, 169, 168), idx(169, 173, 174), idx(174, 170, 169), idx(170, 174, 175), idx(175, 171, 170), 
		idx(111, 115, 176), idx(176, 172, 111), idx(172, 176, 177), idx(177, 173, 172), idx(173, 177, 178), idx(178, 174, 173), idx(174, 178, 179), idx(179, 175, 174), idx(115, 119, 180), idx(180, 176, 115), 
		idx(176, 180, 181), idx(181, 177, 176), idx(177, 181, 182), idx(182, 178, 177), idx(178, 182, 183), idx(183, 179, 178), idx(119, 123, 184), idx(184, 180, 119), idx(180, 184, 185), idx(185, 181, 180), 
		idx(181, 185, 186), idx(186, 182, 181), idx(182, 186, 187), idx(187, 183, 182), idx(123, 127, 188), idx(188, 184, 123), idx(184, 188, 189), idx(189, 185, 184), idx(185, 189, 190), idx(190, 186, 185), 
		idx(186, 190, 191), idx(191, 187, 186), idx(127, 131, 192), idx(192, 188, 127), idx(188, 192, 193), idx(193, 189, 188), idx(189, 193, 194), idx(194, 190, 189), idx(190, 194, 195), idx(195, 191, 190), 
		idx(131, 135, 196), idx(196, 192, 131), idx(192, 196, 197), idx(197, 193, 192), idx(193, 197, 198), idx(198, 194, 193), idx(194, 198, 199), idx(199, 195, 194), idx(135, 139, 200), idx(200, 196, 135), 
		idx(196, 200, 201), idx(201, 197, 196), idx(197, 201, 202), idx(202, 198, 197), idx(198, 202, 203), idx(203, 199, 198), idx(139, 143, 204), idx(204, 200, 139), idx(200, 204, 205), idx(205, 201, 200), 
		idx(201, 205, 206), idx(206, 202, 201), idx(202, 206, 207), idx(207, 203, 202), idx(143, 87, 145), idx(145, 204, 143), idx(204, 145, 147), idx(147, 205, 204), idx(205, 147, 149), idx(149, 206, 205), 
		idx(206, 149, 151), idx(151, 207, 206), idx(151, 150, 208), idx(208, 209, 151), idx(209, 208, 210), idx(210, 211, 209), idx(211, 210, 212), idx(212, 213, 211), idx(213, 212, 214), idx(214, 214, 213), 
		idx(150, 155, 215), idx(215, 208, 150), idx(208, 215, 216), idx(216, 210, 208), idx(210, 216, 217), idx(217, 212, 210), idx(212, 217, 214), idx(214, 214, 212), idx(155, 159, 218), idx(218, 215, 155), 
		idx(215, 218, 219), idx(219, 216, 215), idx(216, 219, 220), idx(220, 217, 216), idx(217, 220, 214), idx(214, 214, 217), idx(159, 163, 221), idx(221, 218, 159), idx(218, 221, 222), idx(222, 219, 218), 
		idx(219, 222, 223), idx(223, 220, 219), idx(220, 223, 214), idx(214, 214, 220), idx(163, 167, 224), idx(224, 221, 163), idx(221, 224, 225), idx(225, 222, 221), idx(222, 225, 226), idx(226, 223, 222), 
		idx(223, 226, 214), idx(214, 214, 223), idx(167, 171, 227), idx(227, 224, 167), idx(224, 227, 228), idx(228, 225, 224), idx(225, 228, 229), idx(229, 226, 225), idx(226, 229, 214), idx(214, 214, 226), 
		idx(171, 175, 230), idx(230, 227, 171), idx(227, 230, 231), idx(231, 228, 227), idx(228, 231, 232), idx(232, 229, 228), idx(229, 232, 214), idx(214, 214, 229), idx(175, 179, 233), idx(233, 230, 175), 
		idx(230, 233, 234), idx(234, 231, 230), idx(231, 234, 235), idx(235, 232, 231), idx(232, 235, 214), idx(214, 214, 232), idx(179, 183, 236), idx(236, 233, 179), idx(233, 236, 237), idx(237, 234, 233), 
		idx(234, 237, 238), idx(238, 235, 234), idx(235, 238, 214), idx(214, 214, 235), idx(183, 187, 239), idx(239, 236, 183), idx(236, 239, 240), idx(240, 237, 236), idx(237, 240, 241), idx(241, 238, 237), 
		idx(238, 241, 214), idx(214, 214, 238), idx(187, 191, 242), idx(242, 239, 187), idx(239, 242, 243), idx(243, 240, 239), idx(240, 243, 244), idx(244, 241, 240), idx(241, 244, 214), idx(214, 214, 241), 
		idx(191, 195, 245), idx(245, 242, 191), idx(242, 245, 246), idx(246, 243, 242), idx(243, 246, 247), idx(247, 244, 243), idx(244, 247, 214), idx(214, 214, 244), idx(195, 199, 248), idx(248, 245, 195), 
		idx(245, 248, 249), idx(249, 246, 245), idx(246, 249, 250), idx(250, 247, 246), idx(247, 250, 214), idx(214, 214, 247), idx(199, 203, 251), idx(251, 248, 199), idx(248, 251, 252), idx(252, 249, 248), 
		idx(249, 252, 253), idx(253, 250, 249), idx(250, 253, 214), idx(214, 214, 250), idx(203, 207, 254), idx(254, 251, 203), idx(251, 254, 255), idx(255, 252, 251), idx(252, 255, 256), idx(256, 253, 252), 
		idx(253, 256, 214), idx(214, 214, 253), idx(207, 151, 209), idx(209, 254, 207), idx(254, 209, 211), idx(211, 255, 254), idx(255, 211, 213), idx(213, 256, 255), idx(256, 213, 214), idx(214, 214, 256), 
		idx(257, 258, 259), idx(259, 260, 257), idx(260, 259, 261), idx(261, 262, 260), idx(262, 261, 263), idx(263, 264, 262), idx(264, 263, 265), idx(265, 266, 264), idx(258, 267, 268), idx(268, 259, 258), 
		idx(259, 268, 269), idx(269, 261, 259), idx(261, 269, 270), idx(270, 263, 261), idx(263, 270, 271), idx(271, 265, 263), idx(267, 272, 273), idx(273, 268, 267), idx(268, 273, 274), idx(274, 269, 268), 
		idx(269, 274, 275), idx(275, 270, 269), idx(270, 275, 276), idx(276, 271, 270), idx(272, 277, 278), idx(278, 273, 272), idx(273, 278, 279), idx(279, 274, 273), idx(274, 279, 280), idx(280, 275, 274), 
		idx(275, 280, 281), idx(281, 276, 275), idx(277, 282, 283), idx(283, 278, 277), idx(278, 283, 284), idx(284, 279, 278), idx(279, 284, 285), idx(285, 280, 279), idx(280, 285, 286), idx(286, 281, 280), 
		idx(282, 287, 288), idx(288, 283, 282), idx(283, 288, 289), idx(289, 284, 283), idx(284, 289, 290), idx(290, 285, 284), idx(285, 290, 291), idx(291, 286, 285), idx(287, 292, 293), idx(293, 288, 287), 
		idx(288, 293, 294), idx(294, 289, 288), idx(289, 294, 295), idx(295, 290, 289), idx(290, 295, 296), idx(296, 291, 290), idx(292, 257, 260), idx(260, 293, 292), idx(293, 260, 262), idx(262, 294, 293), 
		idx(294, 262, 264), idx(264, 295, 294), idx(295, 264, 266), idx(266, 296, 295), idx(266, 265, 297), idx(297, 298, 266), idx(298, 297, 299), idx(299, 300, 298), idx(300, 299, 301), idx(301, 302, 300), 
		idx(302, 301, 303), idx(303, 115, 302), idx(265, 271, 304), idx(304, 297, 265), idx(297, 304, 305), idx(305, 299, 297), idx(299, 305, 306), idx(306, 301, 299), idx(301, 306, 307), idx(307, 303, 301), 
		idx(271, 276, 308), idx(308, 304, 271), idx(304, 308, 309), idx(309, 305, 304), idx(305, 309, 310), idx(310, 306, 305), idx(306, 310, 311), idx(311, 307, 306), idx(276, 281, 312), idx(312, 308, 276), 
		idx(308, 312, 313), idx(313, 309, 308), idx(309, 313, 314), idx(314, 310, 309), idx(310, 314, 315), idx(315, 311, 310), idx(281, 286, 316), idx(316, 312, 281), idx(312, 316, 317), idx(317, 313, 312), 
		idx(313, 317, 318), idx(318, 314, 313), idx(314, 318, 319), idx(319, 315, 314), idx(286, 291, 320), idx(320, 316, 286), idx(316, 320, 321), idx(321, 317, 316), idx(317, 321, 322), idx(322, 318, 317), 
		idx(318, 322, 323), idx(323, 319, 318), idx(291, 296, 324), idx(324, 320, 291), idx(320, 324, 325), idx(325, 321, 320), idx(321, 325, 326), idx(326, 322, 321), idx(322, 326, 327), idx(327, 323, 322), 
		idx(296, 266, 298), idx(298, 324, 296), idx(324, 298, 300), idx(300, 325, 324), idx(325, 300, 302), idx(302, 326, 325), idx(326, 302, 115), idx(115, 327, 326), idx(328, 329, 330), idx(330, 331, 328), 
		idx(331, 330, 332), idx(332, 333, 331), idx(333, 332, 334), idx(334, 335, 333), idx(335, 334, 336), idx(336, 337, 335), idx(329, 338, 339), idx(339, 330, 329), idx(330, 339, 340), idx(340, 332, 330), 
		idx(332, 340, 341), idx(341, 334, 332), idx(334, 341, 342), idx(342, 336, 334), idx(338, 343, 344), idx(344, 339, 338), idx(339, 344, 345), idx(345, 340, 339), idx(340, 345, 346), idx(346, 341, 340), 
		idx(341, 346, 347), idx(347, 342, 341), idx(343, 348, 349), idx(349, 344, 343), idx(344, 349, 350), idx(350, 345, 344), idx(345, 350, 351), idx(351, 346, 345), idx(346, 351, 352), idx(352, 347, 346), 
		idx(348, 353, 354), idx(354, 349, 348), idx(349, 354, 355), idx(355, 350, 349), idx(350, 355, 356), idx(356, 351, 350), idx(351, 356, 357), idx(357, 352, 351), idx(353, 358, 359), idx(359, 354, 353), 
		idx(354, 359, 360), idx(360, 355, 354), idx(355, 360, 361), idx(361, 356, 355), idx(356, 361, 362), idx(362, 357, 356), idx(358, 363, 364), idx(364, 359, 358), idx(359, 364, 365), idx(365, 360, 359), 
		idx(360, 365, 366), idx(366, 361, 360), idx(361, 366, 367), idx(367, 362, 361), idx(363, 328, 331), idx(331, 364, 363), idx(364, 331, 333), idx(333, 365, 364), idx(365, 333, 335), idx(335, 366, 365), 
		idx(366, 335, 337), idx(337, 367, 366), idx(337, 336, 368), idx(368, 369, 337), idx(369, 368, 370), idx(370, 371, 369), idx(371, 370, 372), idx(372, 373, 371), idx(373, 372, 374), idx(374, 375, 373), 
		idx(336, 342, 376), idx(376, 368, 336), idx(368, 376, 377), idx(377, 370, 368), idx(370, 377, 378), idx(378, 372, 370), idx(372, 378, 379), idx(379, 374, 372), idx(342, 347, 380), idx(380, 376, 342), 
		idx(376, 380, 381), idx(381, 377, 376), idx(377, 381, 382), idx(382, 378, 377), idx(378, 382, 383), idx(383, 379, 378), idx(347, 352, 384), idx(384, 380, 347), idx(380, 384, 385), idx(385, 381, 380), 
		idx(381, 385, 386), idx(386, 382, 381), idx(382, 386, 387), idx(387, 383, 382), idx(352, 357, 388), idx(388, 384, 352), idx(384, 388, 389), idx(389, 385, 384), idx(385, 389, 390), idx(390, 386, 385), 
		idx(386, 390, 391), idx(391, 387, 386), idx(357, 362, 392), idx(392, 388, 357), idx(388, 392, 393), idx(393, 389, 388), idx(389, 393, 394), idx(394, 390, 389), idx(390, 394, 395), idx(395, 391, 390), 
		idx(362, 367, 396), idx(396, 392, 362), idx(392, 396, 397), idx(397, 393, 392), idx(393, 397, 398), idx(398, 394, 393), idx(394, 398, 399), idx(399, 395, 394), idx(367, 337, 369), idx(369, 396, 367), 
		idx(396, 369, 371), idx(371, 397, 396), idx(397, 371, 373), idx(373, 398, 397), idx(398, 373, 375), idx(375, 399, 398), idx(400, 400, 401), idx(401, 402, 400), idx(402, 401, 403), idx(403, 404, 402), 
		idx(404, 403, 405), idx(405, 406, 404), idx(406, 405, 407), idx(407, 408, 406), idx(400, 400, 409), idx(409, 401, 400), idx(401, 409, 410), idx(410, 403, 401), idx(403, 410, 411), idx(411, 405, 403), 
		idx(405, 411, 412), idx(412, 407, 405), idx(400, 400, 413), idx(413, 409, 400), idx(409, 413, 414), idx(414, 410, 409), idx(410, 414, 415), idx(415, 411, 410), idx(411, 415, 416), idx(416, 412, 411), 
		idx(400, 400, 417), idx(417, 413, 400), idx(413, 417, 418), idx(418, 414, 413), idx(414, 418, 419), idx(419, 415, 414), idx(415, 419, 420), idx(420, 416, 415), idx(400, 400, 421), idx(421, 417, 400), 
		idx(417, 421, 422), idx(422, 418, 417), idx(418, 422, 423), idx(423, 419, 418), idx(419, 423, 424), idx(424, 420, 419), idx(400, 400, 425), idx(425, 421, 400), idx(421, 425, 426), idx(426, 422, 421), 
		idx(422, 426, 427), idx(427, 423, 422), idx(423, 427, 428), idx(428, 424, 423), idx(400, 400, 429), idx(429, 425, 400), idx(425, 429, 430), idx(430, 426, 425), idx(426, 430, 431), idx(431, 427, 426), 
		idx(427, 431, 432), idx(432, 428, 427), idx(400, 400, 433), idx(433, 429, 400), idx(429, 433, 434), idx(434, 430, 429), idx(430, 434, 435), idx(435, 431, 430), idx(431, 435, 436), idx(436, 432, 431), 
		idx(400, 400, 437), idx(437, 433, 400), idx(433, 437, 438), idx(438, 434, 433), idx(434, 438, 439), idx(439, 435, 434), idx(435, 439, 440), idx(440, 436, 435), idx(400, 400, 441), idx(441, 437, 400), 
		idx(437, 441, 442), idx(442, 438, 437), idx(438, 442, 443), idx(443, 439, 438), idx(439, 443, 444), idx(444, 440, 439), idx(400, 400, 445), idx(445, 441, 400), idx(441, 445, 446), idx(446, 442, 441), 
		idx(442, 446, 447), idx(447, 443, 442), idx(443, 447, 448), idx(448, 444, 443), idx(400, 400, 449), idx(449, 445, 400), idx(445, 449, 450), idx(450, 446, 445), idx(446, 450, 451), idx(451, 447, 446), 
		idx(447, 451, 452), idx(452, 448, 447), idx(400, 400, 453), idx(453, 449, 400), idx(449, 453, 454), idx(454, 450, 449), idx(450, 454, 455), idx(455, 451, 450), idx(451, 455, 456), idx(456, 452, 451), 
		idx(400, 400, 457), idx(457, 453, 400), idx(453, 457, 458), idx(458, 454, 453), idx(454, 458, 459), idx(459, 455, 454), idx(455, 459, 460), idx(460, 456, 455), idx(400, 400, 461), idx(461, 457, 400), 
		idx(457, 461, 462), idx(462, 458, 457), idx(458, 462, 463), idx(463, 459, 458), idx(459, 463, 464), idx(464, 460, 459), idx(400, 400, 402), idx(402, 461, 400), idx(461, 402, 404), idx(404, 462, 461), 
		idx(462, 404, 406), idx(406, 463, 462), idx(463, 406, 408), idx(408, 464, 463), idx(408, 407, 465), idx(465, 466, 408), idx(466, 465, 467), idx(467, 468, 466), idx(468, 467, 469), idx(469, 470, 468), 
		idx(470, 469, 471), idx(471, 472, 470), idx(407, 412, 473), idx(473, 465, 407), idx(465, 473, 474), idx(474, 467, 465), idx(467, 474, 475), idx(475, 469, 467), idx(469, 475, 476), idx(476, 471, 469), 
		idx(412, 416, 477), idx(477, 473, 412), idx(473, 477, 478), idx(478, 474, 473), idx(474, 478, 479), idx(479, 475, 474), idx(475, 479, 480), idx(480, 476, 475), idx(416, 420, 481), idx(481, 477, 416), 
		idx(477, 481, 482), idx(482, 478, 477), idx(478, 482, 483), idx(483, 479, 478), idx(479, 483, 484), idx(484, 480, 479), idx(420, 424, 485), idx(485, 481, 420), idx(481, 485, 486), idx(486, 482, 481), 
		idx(482, 486, 487), idx(487, 483, 482), idx(483, 487, 488), idx(488, 484, 483), idx(424, 428, 489), idx(489, 485, 424), idx(485, 489, 490), idx(490, 486, 485), idx(486, 490, 491), idx(491, 487, 486), 
		idx(487, 491, 492), idx(492, 488, 487), idx(428, 432, 493), idx(493, 489, 428), idx(489, 493, 494), idx(494, 490, 489), idx(490, 494, 495), idx(495, 491, 490), idx(491, 495, 496), idx(496, 492, 491), 
		idx(432, 436, 497), idx(497, 493, 432), idx(493, 497, 498), idx(498, 494, 493), idx(494, 498, 499), idx(499, 495, 494), idx(495, 499, 500), idx(500, 496, 495), idx(436, 440, 501), idx(501, 497, 436), 
		idx(497, 501, 502), idx(502, 498, 497), idx(498, 502, 503), idx(503, 499, 498), idx(499, 503, 504), idx(504, 500, 499), idx(440, 444, 505), idx(505, 501, 440), idx(501, 505, 506), idx(506, 502, 501), 
		idx(502, 506, 507), idx(507, 503, 502), idx(503, 507, 508), idx(508, 504, 503), idx(444, 448, 509), idx(509, 505, 444), idx(505, 509, 510), idx(510, 506, 505), idx(506, 510, 511), idx(511, 507, 506), 
		idx(507, 511, 512), idx(512, 508, 507), idx(448, 452, 513), idx(513, 509, 448), idx(509, 513, 514), idx(514, 510, 509), idx(510, 514, 515), idx(515, 511, 510), idx(511, 515, 516), idx(516, 512, 511), 
		idx(452, 456, 517), idx(517, 513, 452), idx(513, 517, 518), idx(518, 514, 513), idx(514, 518, 519), idx(519, 515, 514), idx(515, 519, 520), idx(520, 516, 515), idx(456, 460, 521), idx(521, 517, 456), 
		idx(517, 521, 522), idx(522, 518, 517), idx(518, 522, 523), idx(523, 519, 518), idx(519, 523, 524), idx(524, 520, 519), idx(460, 464, 525), idx(525, 521, 460), idx(521, 525, 526), idx(526, 522, 521), 
		idx(522, 526, 527), idx(527, 523, 522), idx(523, 527, 528), idx(528, 524, 523), idx(464, 408, 466), idx(466, 525, 464), idx(525, 466, 468), idx(468, 526, 525), idx(526, 468, 470), idx(470, 527, 526), 
		idx(527, 470, 472), idx(472, 528, 527)
	);

end package renderer_mesh;
