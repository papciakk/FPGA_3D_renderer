use work.common.all;

package renderer_mesh is

	--	constant vertices : vertex_arr_t(0 to 4) := (
	--		point2d(18, 83),
	--		point2d(130, 19),
	--		point2d(170, 120),
	--		point2d(40, 115),
	--		point2d(172, 26)
	--	);
	--
	--	constant indices : indices_arr_t(0 to 2) := (
	--		idx(1, 0, 2),
	--		idx(3, 0, 2),
	--		idx(1, 2, 4)
	--	);

	--	constant vertices : vertex_arr_t(0 to 7)  := (
	--		point2d(66, 80),
	--		point2d(32, 81),
	--		point2d(80, 110),
	--		point2d(113, 93),
	--		point2d(74, 31),
	--		point2d(40, 32),
	--		point2d(19, 72),
	--		point2d(120, 69)
	--	);
	--	constant indices  : indices_arr_t := (
	--		idx(0, 5, 4),
	--		idx(1, 6, 5),
	--		idx(7, 3, 4),
	--		idx(1, 5, 0),
	--		idx(0, 4, 3),
	--		idx(0, 3, 2),
	--		idx(1, 0, 2)
	--	);

	constant vertices : vertex_arr_t(0 to 67) := (
	point2d(7, 3),
	point2d(7, 42),
	point2d(12, 42),
	point2d(12, 9),
	point2d(15, 3),
	point2d(24, 31),
	point2d(23, 42),
	point2d(26, 36),
	point2d(28, 42),
	point2d(39, 10),
	point2d(28, 30),
	point2d(37, 3),
	point2d(44, 3),
	point2d(44, 42),
	point2d(39, 42),
	point2d(66, 7),
	point2d(54, 42),
	point2d(58, 30),
	point2d(65, 8),
	point2d(65, 10),
	point2d(65, 11),
	point2d(64, 12),
	point2d(78, 42),
	point2d(84, 42),
	point2d(69, 3),
	point2d(74, 30),
	point2d(63, 3),
	point2d(48, 42),
	point2d(66, 8),
	point2d(66, 9),
	point2d(67, 10),
	point2d(67, 12),
	point2d(67, 13),
	point2d(64, 14),
	point2d(64, 13),
	point2d(63, 15),
	point2d(59, 26),
	point2d(72, 26),
	point2d(68, 15),
	point2d(68, 14),
	point2d(99, 22),
	point2d(84, 42),
	point2d(90, 42),
	point2d(100, 29),
	point2d(102, 26),
	point2d(105, 22),
	point2d(118, 3),
	point2d(113, 3),
	point2d(105, 14),
	point2d(105, 14),
	point2d(104, 15),
	point2d(104, 15),
	point2d(103, 16),
	point2d(103, 17),
	point2d(113, 42),
	point2d(120, 42),
	point2d(104, 28),
	point2d(92, 3),
	point2d(86, 3),
	point2d(99, 13),
	point2d(100, 14),
	point2d(100, 15),
	point2d(101, 16),
	point2d(101, 16),
	point2d(102, 17),
	point2d(103, 17),
	point2d(102, 17),
	point2d(102, 18)
);
constant indices : indices_arr_t(0 to 63) := (
	idx(0, 1, 2),
	idx(0, 2, 3),
	idx(4, 0, 3),
	idx(5, 4, 3),
	idx(5, 3, 6),
	idx(7, 5, 6),
	idx(7, 6, 8),
	idx(7, 8, 9),
	idx(10, 7, 9),
	idx(11, 10, 9),
	idx(12, 11, 9),
	idx(13, 12, 9),
	idx(13, 9, 14),
	idx(15, 16, 17),
	idx(18, 15, 17),
	idx(19, 18, 17),
	idx(20, 19, 17),
	idx(21, 20, 17),
	idx(22, 23, 24),
	idx(25, 22, 24),
	idx(26, 27, 16),
	idx(26, 16, 15),
	idx(24, 26, 15),
	idx(25, 24, 15),
	idx(25, 15, 28),
	idx(25, 28, 29),
	idx(25, 29, 30),
	idx(25, 30, 31),
	idx(25, 31, 32),
	idx(33, 34, 21),
	idx(35, 33, 21),
	idx(36, 35, 21),
	idx(36, 21, 17),
	idx(36, 17, 25),
	idx(37, 36, 25),
	idx(38, 37, 25),
	idx(38, 25, 32),
	idx(39, 38, 32),
	idx(40, 41, 42),
	idx(40, 42, 43),
	idx(40, 43, 44),
	idx(45, 46, 47),
	idx(45, 47, 48),
	idx(45, 48, 49),
	idx(45, 49, 50),
	idx(45, 50, 51),
	idx(45, 51, 52),
	idx(45, 52, 53),
	idx(54, 55, 45),
	idx(56, 54, 45),
	idx(44, 56, 45),
	idx(57, 58, 40),
	idx(59, 57, 40),
	idx(60, 59, 40),
	idx(61, 60, 40),
	idx(62, 61, 40),
	idx(63, 62, 40),
	idx(64, 63, 40),
	idx(45, 53, 65),
	idx(66, 64, 40),
	idx(67, 66, 40),
	idx(45, 65, 67),
	idx(40, 44, 45),
	idx(67, 40, 45)
);
end package renderer_mesh;
