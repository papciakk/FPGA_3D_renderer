library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity triangle_renderer is
	port(
		clk : in std_logic;
		rst : in std_logic
	);
end entity triangle_renderer;

architecture bahavioral of triangle_renderer is
	
begin

end architecture bahavioral;
