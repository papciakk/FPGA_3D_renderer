use work.common.all;

package renderer_mesh is
	constant vertices : vertex_attr_arr_t(0 to 137) := (
		va(10059, -2420, 4953, 0, 124, 130), va(7156, -8209, 824, 37, 197, 182), va(7173, -8632, 1389, 114, 63, 236), va(10086, -2826, 5529, 109, 53, 229), va(7666, -8621, 526, 202, 25, 139), va(10776, -2420, 4953, 233, 86, 183), va(43, -10575, -862, 126, 228, 203), va(43, -10998, -303, 126, 68, 239), va(43, -11155, -1280, 127, 0, 121), va(-7308, -8209, 824, 219, 208, 157), va(-7113, -8632, 1389, 137, 77, 243), 
		va(-7574, -8621, 526, 51, 25, 138), va(-9973, -2420, 4953, 253, 123, 129), va(-9994, -2826, 5529, 145, 52, 228), va(-10689, -2420, 4953, 20, 87, 183), va(-7070, 3369, 9083, 216, 51, 78), va(-7080, 2973, 9663, 139, 43, 222), va(-7574, 3787, 9376, 51, 148, 226), va(43, 5735, 10770, 127, 21, 56), va(43, 5344, 11356, 127, 39, 218), va(43, 6321, 11188, 127, 173, 245), 
		va(7156, 3369, 9083, 37, 51, 78), va(7173, 2973, 9663, 114, 43, 222), va(7666, 3787, 9376, 202, 148, 226), va(9414, -6809, -5019, 212, 34, 108), va(13239, 813, 417, 248, 104, 158), va(10206, -4454, -9685, 216, 62, 63), va(14357, 3814, -3787, 253, 135, 115), va(43, -9924, -7238, 127, 6, 87), va(43, -7835, -12094, 127, 32, 42), va(-9321, -6809, -5019, 41, 34, 108), 
		va(-10114, -4454, -9685, 37, 62, 63), va(-13147, 813, 417, 5, 104, 158), va(-14265, 3814, -3787, 0, 135, 115), va(-9321, 8442, 5860, 41, 174, 208), va(-10114, 12089, 2116, 37, 207, 167), va(43, 11557, 8079, 127, 203, 228), va(43, 15464, 4525, 127, 237, 188), va(9414, 8442, 5860, 212, 174, 208), va(10206, 12089, 2116, 216, 207, 167), va(8936, -1280, -11953, 200, 109, 24), 
		va(12566, 5957, -6787, 231, 169, 67), va(7666, 727, -12577, 179, 143, 12), va(10776, 6929, -8155, 201, 186, 43), va(43, -4237, -14058, 127, 84, 7), va(43, -1806, -14384, 127, 125, 0), va(-8844, -1280, -11953, 53, 109, 24), va(-7574, 727, -12577, 74, 143, 12), va(-12474, 5957, -6787, 22, 169, 67), va(-10689, 6929, -8155, 52, 186, 43), va(-8844, 13196, -1627, 53, 229, 110), 
		va(-7574, 13136, -3727, 74, 229, 74), va(43, 16153, 482, 127, 253, 128), va(43, 15670, -1920, 127, 247, 86), va(8936, 13196, -1627, 200, 229, 110), va(7666, 13136, -3727, 179, 229, 74), va(6570, 2045, -12544, 152, 176, 13), va(9235, 7357, -8752, 163, 197, 27), va(43, 7553, -9028, 127, 200, 23), va(43, -124, -14091, 127, 168, 6), va(-6478, 2045, -12544, 101, 176, 13), 
		va(-9142, 7357, -8752, 90, 197, 27), va(-6478, 12669, -4964, 101, 218, 42), va(43, 14840, -3418, 127, 227, 48), va(6570, 12669, -4964, 152, 218, 42), va(-11405, -857, 2767, 131, 201, 23), va(-11047, -2637, 2490, 124, 7, 84), va(-17976, -2463, 2240, 124, 10, 75), va(-17216, -743, 2604, 162, 199, 28), va(-20347, -1237, 520, 89, 19, 70), va(-19273, 75, 1459, 245, 157, 92), 
		va(-10689, -1796, 4080, 120, 53, 230), va(-18736, -1562, 3749, 70, 59, 218), va(-21421, 75, 1459, 1, 113, 143), va(-11047, -16, 4357, 124, 206, 225), va(-17976, 157, 4112, 125, 215, 218), va(-20347, 1383, 2392, 92, 218, 208), va(-18806, 1030, -2658, 111, 32, 43), va(-18112, 1942, -1161, 230, 85, 187), va(-13906, 3125, -5594, 84, 82, 16), va(-14265, 3814, -3787, 205, 72, 210), 
		va(-19495, 2745, -2284, 28, 172, 61), va(-13548, 5062, -5534, 54, 186, 41), va(-18806, 3657, -786, 113, 235, 190), va(-13906, 5746, -3722, 88, 247, 137), va(12208, 1633, -727, 65, 63, 217), va(12208, 461, -5187, 168, 50, 34), va(18198, -1172, -998, 147, 23, 56), va(17129, 75, 1459, 38, 71, 199), va(21508, -3510, 4172, 126, 3, 98), va(19365, -2420, 4953, 35, 70, 194), 
		va(12208, 5062, -5534, 210, 183, 48), va(19273, 1557, -618, 224, 176, 62), va(23657, -2420, 4953, 209, 187, 51), va(12208, 6229, -1074, 170, 238, 169), va(18198, 2805, 1839, 150, 228, 200), va(21508, -1323, 5729, 133, 201, 229), va(22414, -3570, 4720, 156, 9, 164), va(20260, -2653, 5279, 132, 46, 224), va(21508, -3071, 4487, 167, 228, 192), va(20081, -2420, 4953, 241, 157, 81), 
		va(24574, -2740, 5404, 248, 108, 160), va(22941, -2420, 4953, 86, 57, 225), va(22414, -1823, 5963, 173, 133, 245), va(21508, -1763, 5420, 170, 39, 46), va(43, -5534, 9321, 127, 53, 230), va(1698, -6180, 7379, 213, 35, 106), va(2371, -4834, 8339, 248, 105, 156), va(1063, -4492, 6109, 202, 25, 138), va(1475, -3662, 6701, 234, 87, 182), va(43, -6728, 6988, 126, 6, 86), 
		va(43, -4829, 5870, 126, 0, 120), va(-1606, -6180, 7379, 40, 35, 106), va(-971, -4492, 6109, 51, 25, 138), va(-2278, -4834, 8339, 5, 105, 156), va(-1383, -3662, 6701, 19, 87, 182), va(-1606, -3488, 9300, 40, 175, 206), va(-971, -2837, 7292, 51, 148, 226), va(43, -2940, 9690, 127, 204, 227), va(43, -2501, 7531, 127, 174, 244), va(1698, -3488, 9300, 213, 175, 206), 
		va(1063, -2837, 7292, 202, 148, 226), va(4237, -6451, 3391, 151, 36, 212), va(5946, -3044, 5827, 161, 56, 226), va(6646, -7797, 1117, 153, 34, 209), va(9349, -2420, 4953, 165, 56, 225), va(43, -7846, 2398, 127, 27, 206), va(43, -9989, -450, 127, 25, 203), va(-4145, -6451, 3391, 102, 36, 212), va(-6560, -7797, 1117, 100, 34, 209), va(-5860, -3044, 5827, 92, 56, 226), 
		va(-9256, -2420, 4953, 88, 56, 225), va(-4145, 368, 8258, 102, 76, 240), va(-6560, 2957, 8790, 100, 78, 241), va(43, 1763, 9256, 127, 84, 246), va(43, 5154, 10352, 127, 87, 247), va(4237, 368, 8258, 151, 76, 240), va(6646, 2957, 8790, 153, 78, 241)
	);

	constant indices : indices_arr_t(0 to 255) := (
		idx(0, 1, 2), idx(2, 3, 0), 
		idx(3, 2, 4), idx(4, 5, 3), idx(1, 6, 7), idx(7, 2, 1), idx(2, 7, 8), idx(8, 4, 2), idx(6, 9, 10), idx(10, 7, 6), idx(7, 10, 11), idx(11, 8, 7), 
		idx(9, 12, 13), idx(13, 10, 9), idx(10, 13, 14), idx(14, 11, 10), idx(12, 15, 16), idx(16, 13, 12), idx(13, 16, 17), idx(17, 14, 13), idx(15, 18, 19), idx(19, 16, 15), 
		idx(16, 19, 20), idx(20, 17, 16), idx(18, 21, 22), idx(22, 19, 18), idx(19, 22, 23), idx(23, 20, 19), idx(21, 0, 3), idx(3, 22, 21), idx(22, 3, 5), idx(5, 23, 22), 
		idx(5, 4, 24), idx(24, 25, 5), idx(25, 24, 26), idx(26, 27, 25), idx(4, 8, 28), idx(28, 24, 4), idx(24, 28, 29), idx(29, 26, 24), idx(8, 11, 30), idx(30, 28, 8), 
		idx(28, 30, 31), idx(31, 29, 28), idx(11, 14, 32), idx(32, 30, 11), idx(30, 32, 33), idx(33, 31, 30), idx(14, 17, 34), idx(34, 32, 14), idx(32, 34, 35), idx(35, 33, 32), 
		idx(17, 20, 36), idx(36, 34, 17), idx(34, 36, 37), idx(37, 35, 34), idx(20, 23, 38), idx(38, 36, 20), idx(36, 38, 39), idx(39, 37, 36), idx(23, 5, 25), idx(25, 38, 23), 
		idx(38, 25, 27), idx(27, 39, 38), idx(27, 26, 40), idx(40, 41, 27), idx(41, 40, 42), idx(42, 43, 41), idx(26, 29, 44), idx(44, 40, 26), idx(40, 44, 45), idx(45, 42, 40), 
		idx(29, 31, 46), idx(46, 44, 29), idx(44, 46, 47), idx(47, 45, 44), idx(31, 33, 48), idx(48, 46, 31), idx(46, 48, 49), idx(49, 47, 46), idx(33, 35, 50), idx(50, 48, 33), 
		idx(48, 50, 51), idx(51, 49, 48), idx(35, 37, 52), idx(52, 50, 35), idx(50, 52, 53), idx(53, 51, 50), idx(37, 39, 54), idx(54, 52, 37), idx(52, 54, 55), idx(55, 53, 52), 
		idx(39, 27, 41), idx(41, 54, 39), idx(54, 41, 43), idx(43, 55, 54), idx(43, 42, 56), idx(56, 57, 43), idx(57, 56, 58), idx(58, 58, 57), idx(42, 45, 59), idx(59, 56, 42), 
		idx(56, 59, 58), idx(58, 58, 56), idx(45, 47, 60), idx(60, 59, 45), idx(59, 60, 58), idx(58, 58, 59), idx(47, 49, 61), idx(61, 60, 47), idx(60, 61, 58), idx(58, 58, 60), 
		idx(49, 51, 62), idx(62, 61, 49), idx(61, 62, 58), idx(58, 58, 61), idx(51, 53, 63), idx(63, 62, 51), idx(62, 63, 58), idx(58, 58, 62), idx(53, 55, 64), idx(64, 63, 53), 
		idx(63, 64, 58), idx(58, 58, 63), idx(55, 43, 57), idx(57, 64, 55), idx(64, 57, 58), idx(58, 58, 64), idx(65, 66, 67), idx(67, 68, 65), idx(68, 67, 69), idx(69, 70, 68), 
		idx(66, 71, 72), idx(72, 67, 66), idx(67, 72, 73), idx(73, 69, 67), idx(71, 74, 75), idx(75, 72, 71), idx(72, 75, 76), idx(76, 73, 72), idx(74, 65, 68), idx(68, 75, 74), 
		idx(75, 68, 70), idx(70, 76, 75), idx(70, 69, 77), idx(77, 78, 70), idx(78, 77, 79), idx(79, 80, 78), idx(69, 73, 81), idx(81, 77, 69), idx(77, 81, 82), idx(82, 79, 77), 
		idx(73, 76, 83), idx(83, 81, 73), idx(81, 83, 84), idx(84, 82, 81), idx(76, 70, 78), idx(78, 83, 76), idx(83, 78, 80), idx(80, 84, 83), idx(85, 86, 87), idx(87, 88, 85), 
		idx(88, 87, 89), idx(89, 90, 88), idx(86, 91, 92), idx(92, 87, 86), idx(87, 92, 93), idx(93, 89, 87), idx(91, 94, 95), idx(95, 92, 91), idx(92, 95, 96), idx(96, 93, 92), 
		idx(94, 85, 88), idx(88, 95, 94), idx(95, 88, 90), idx(90, 96, 95), idx(90, 89, 97), idx(97, 98, 90), idx(98, 97, 99), idx(99, 100, 98), idx(89, 93, 101), idx(101, 97, 89), 
		idx(97, 101, 102), idx(102, 99, 97), idx(93, 96, 103), idx(103, 101, 93), idx(101, 103, 104), idx(104, 102, 101), idx(96, 90, 98), idx(98, 103, 96), idx(103, 98, 100), idx(100, 104, 103), 
		idx(105, 105, 106), idx(106, 107, 105), idx(107, 106, 108), idx(108, 109, 107), idx(105, 105, 110), idx(110, 106, 105), idx(106, 110, 111), idx(111, 108, 106), idx(105, 105, 112), idx(112, 110, 105), 
		idx(110, 112, 113), idx(113, 111, 110), idx(105, 105, 114), idx(114, 112, 105), idx(112, 114, 115), idx(115, 113, 112), idx(105, 105, 116), idx(116, 114, 105), idx(114, 116, 117), idx(117, 115, 114), 
		idx(105, 105, 118), idx(118, 116, 105), idx(116, 118, 119), idx(119, 117, 116), idx(105, 105, 120), idx(120, 118, 105), idx(118, 120, 121), idx(121, 119, 118), idx(105, 105, 107), idx(107, 120, 105), 
		idx(120, 107, 109), idx(109, 121, 120), idx(109, 108, 122), idx(122, 123, 109), idx(123, 122, 124), idx(124, 125, 123), idx(108, 111, 126), idx(126, 122, 108), idx(122, 126, 127), idx(127, 124, 122), 
		idx(111, 113, 128), idx(128, 126, 111), idx(126, 128, 129), idx(129, 127, 126), idx(113, 115, 130), idx(130, 128, 113), idx(128, 130, 131), idx(131, 129, 128), idx(115, 117, 132), idx(132, 130, 115), 
		idx(130, 132, 133), idx(133, 131, 130), idx(117, 119, 134), idx(134, 132, 117), idx(132, 134, 135), idx(135, 133, 132), idx(119, 121, 136), idx(136, 134, 119), idx(134, 136, 137), idx(137, 135, 134), 
		idx(121, 109, 123), idx(123, 136, 121), idx(136, 123, 125), idx(125, 137, 136)
	);

end package renderer_mesh;
