library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.common.all;

entity tile_buffer is

	port 
	(
		clk		: in std_logic;
		addr	: in natural range 0 to 2**16;
		q		: out color_t
	);

end entity;

architecture rtl of tile_buffer is

	type color_buffer_t is array (0 to TILE_RES_X*TILE_RES_Y-1) of color_t;
	signal rom : color_buffer_t := 
	(
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"75", X"75", X"75"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"59", X"59", X"59"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"93", X"93", X"93"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"3B", X"3B", X"3B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"B2", X"B2", X"B2"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FA", X"FA", X"FA"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"D0", X"D0", X"D0"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F0", X"F0", X"F0"), (X"0E", X"0E", X"0E"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"EA", X"EA", X"EA"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"E0", X"E0", X"E0"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"17", X"17", X"17"), (X"F5", X"F5", X"F5"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"C1", X"C1", X"C1"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2B", X"2B", X"2B"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"A3", X"A3", X"A3"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"85", X"85", X"85"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"75", X"75", X"75"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"59", X"59", X"59"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"93", X"93", X"93"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"3B", X"3B", X"3B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"B2", X"B2", X"B2"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FA", X"FA", X"FA"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"D0", X"D0", X"D0"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F0", X"F0", X"F0"), (X"0E", X"0E", X"0E"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"EA", X"EA", X"EA"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"E0", X"E0", X"E0"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"17", X"17", X"17"), (X"F5", X"F5", X"F5"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"C1", X"C1", X"C1"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2B", X"2B", X"2B"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"A3", X"A3", X"A3"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"85", X"85", X"85"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"75", X"75", X"75"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"59", X"59", X"59"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"93", X"93", X"93"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"3B", X"3B", X"3B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"B2", X"B2", X"B2"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FA", X"FA", X"FA"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"D0", X"D0", X"D0"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F0", X"F0", X"F0"), (X"0E", X"0E", X"0E"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"EA", X"EA", X"EA"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"E0", X"E0", X"E0"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"17", X"17", X"17"), (X"F5", X"F5", X"F5"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"C1", X"C1", X"C1"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2B", X"2B", X"2B"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"A3", X"A3", X"A3"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"85", X"85", X"85"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"F4", X"F4", X"F4"), (X"F4", X"F4", X"F4"), (X"F4", X"F4", X"F4"), (X"F4", X"F4", X"F4"), (X"F4", X"F4", X"F4"), (X"F4", X"F4", X"F4"), (X"F8", X"F8", X"F8"), (X"C1", X"C1", X"C1"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"C0", X"C0", X"C0"), (X"FC", X"FC", X"FC"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FD", X"FD", X"FD"), (X"B3", X"B3", X"B3"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"CE", X"CE", X"CE"), (X"FB", X"FB", X"FB"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FD", X"FD", X"FD"), (X"A5", X"A5", X"A5"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"DB", X"DB", X"DB"), (X"FB", X"FB", X"FB"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FB", X"FB", X"FB"), (X"9A", X"9A", X"9A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"E9", X"E9", X"E9"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"F7", X"F7", X"F7"), (X"90", X"90", X"90"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"F0", X"F0", X"F0"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"95", X"95", X"95"), (X"F9", X"F9", X"F9"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FB", X"FB", X"FB"), (X"E3", X"E3", X"E3"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"9E", X"9E", X"9E"), (X"FD", X"FD", X"FD"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FB", X"FB", X"FB"), (X"D5", X"D5", X"D5"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"AC", X"AC", X"AC"), (X"FD", X"FD", X"FD"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FA", X"FA", X"FA"), (X"FC", X"FC", X"FC"), (X"C7", X"C7", X"C7"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"8A", X"8A", X"8A"), (X"B9", X"B9", X"B9"), (X"F9", X"F9", X"F9"), (X"F4", X"F4", X"F4"), (X"F4", X"F4", X"F4"), (X"F4", X"F4", X"F4"), (X"F4", X"F4", X"F4"), (X"F4", X"F4", X"F4"), (X"F4", X"F4", X"F4"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B8", X"B8", X"B8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B7", X"B7", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E1", X"E1", X"E1"), (X"86", X"86", X"86"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E6", X"E6", X"E6"), (X"81", X"81", X"81"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7C", X"7C", X"7C"), (X"E9", X"E9", X"E9"), (X"7C", X"7C", X"7C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"81", X"81", X"81"), (X"E6", X"E6", X"E6"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"BF", X"BF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B0", X"B0", X"B0"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B8", X"B8", X"B8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B7", X"B7", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E1", X"E1", X"E1"), (X"86", X"86", X"86"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E6", X"E6", X"E6"), (X"81", X"81", X"81"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7C", X"7C", X"7C"), (X"E9", X"E9", X"E9"), (X"7C", X"7C", X"7C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"81", X"81", X"81"), (X"E6", X"E6", X"E6"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"BF", X"BF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B0", X"B0", X"B0"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B8", X"B8", X"B8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B7", X"B7", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E1", X"E1", X"E1"), (X"86", X"86", X"86"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E6", X"E6", X"E6"), (X"81", X"81", X"81"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7C", X"7C", X"7C"), (X"E9", X"E9", X"E9"), (X"7C", X"7C", X"7C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"81", X"81", X"81"), (X"E6", X"E6", X"E6"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"BF", X"BF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B0", X"B0", X"B0"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B8", X"B8", X"B8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B7", X"B7", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E1", X"E1", X"E1"), (X"86", X"86", X"86"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E6", X"E6", X"E6"), (X"81", X"81", X"81"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7C", X"7C", X"7C"), (X"E9", X"E9", X"E9"), (X"7C", X"7C", X"7C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"81", X"81", X"81"), (X"E6", X"E6", X"E6"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"BF", X"BF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B0", X"B0", X"B0"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B8", X"B8", X"B8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B7", X"B7", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E1", X"E1", X"E1"), (X"86", X"86", X"86"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E6", X"E6", X"E6"), (X"81", X"81", X"81"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7C", X"7C", X"7C"), (X"E9", X"E9", X"E9"), (X"7C", X"7C", X"7C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"81", X"81", X"81"), (X"E6", X"E6", X"E6"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"BF", X"BF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B0", X"B0", X"B0"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B1", X"BC", X"B8"), (X"6D", X"81", X"7A"), (X"6D", X"81", X"7A"), (X"6D", X"81", X"7A"), (X"6D", X"81", X"7A"), (X"6D", X"81", X"7A"), (X"6D", X"81", X"7A"), (X"6D", X"81", X"7A"), (X"6D", X"81", X"7A"), (X"6D", X"81", X"7A"), (X"B0", X"BB", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E1", X"E1", X"E1"), (X"86", X"86", X"86"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"80", X"80", X"80"), (X"87", X"87", X"87"), (X"A3", X"A3", X"A3"), (X"A7", X"A7", X"A7"), (X"C6", X"C6", X"C6"), (X"F4", X"F4", X"F4"), (X"CD", X"CD", X"CD"), (X"E8", X"E8", X"E8"), (X"E9", X"E9", X"E9"), (X"E9", X"E9", X"E9"), (X"E9", X"E9", X"E9"), (X"E9", X"E9", X"E9"), (X"E9", X"E9", X"E9"), (X"E9", X"E9", X"E9"), (X"E9", X"E9", X"E9"), (X"CD", X"CD", X"CD"), (X"F6", X"F6", X"F6"), (X"C7", X"C7", X"C7"), (X"A9", X"A9", X"A9"), (X"A3", X"A3", X"A3"), (X"89", X"89", X"89"), (X"80", X"80", X"80"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"81", X"81", X"81"), (X"E6", X"E6", X"E6"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"C2", X"B4"), (X"7A", X"7F", X"63"), (X"7A", X"7F", X"63"), (X"7A", X"7F", X"63"), (X"7A", X"7F", X"63"), (X"7A", X"7F", X"63"), (X"7A", X"7F", X"63"), (X"7A", X"7F", X"63"), (X"7A", X"7F", X"63"), (X"7A", X"7F", X"63"), (X"B0", X"B3", X"A2"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E1", X"E1", X"E1"), (X"87", X"87", X"87"), (X"96", X"96", X"96"), (X"B2", X"B2", X"B2"), (X"CB", X"CB", X"CB"), (X"E3", X"E3", X"E3"), (X"FB", X"FB", X"FB"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FD", X"FD", X"FD"), (X"E3", X"E3", X"E3"), (X"CD", X"CD", X"CD"), (X"B4", X"B4", X"B4"), (X"98", X"98", X"98"), (X"82", X"82", X"82"), (X"E6", X"E6", X"E6"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B9", X"B8", X"B8"), (X"7C", X"79", X"7A"), (X"7C", X"79", X"7A"), (X"7C", X"79", X"7A"), (X"7C", X"79", X"7A"), (X"7C", X"79", X"7A"), (X"7C", X"79", X"7A"), (X"7C", X"79", X"7A"), (X"7C", X"79", X"7A"), (X"7C", X"79", X"7A"), (X"B8", X"B7", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8F", X"8F", X"8F"), (X"B4", X"B4", X"B4"), (X"F3", X"F3", X"F3"), (X"FD", X"FD", X"FD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FD", X"FD", X"FD"), (X"F7", X"F7", X"F7"), (X"B6", X"B6", X"B6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"BF", X"C1"), (X"7A", X"79", X"7D"), (X"7A", X"79", X"7D"), (X"7A", X"79", X"7D"), (X"7A", X"79", X"7D"), (X"7A", X"79", X"7D"), (X"7A", X"79", X"7D"), (X"7A", X"79", X"7D"), (X"7A", X"79", X"7D"), (X"7A", X"79", X"7D"), (X"B0", X"AF", X"B1"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"94", X"94", X"94"), (X"C1", X"C1", X"C1"), (X"EB", X"EB", X"EB"), (X"FD", X"FD", X"FD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FE", X"FE", X"FE"), (X"ED", X"ED", X"ED"), (X"C4", X"C4", X"C4"), (X"98", X"98", X"98"), (X"7B", X"7B", X"7B"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"87", X"87", X"87"), (X"B8", X"B8", X"B8"), (X"E7", X"E7", X"E7"), (X"FE", X"FE", X"FE"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FE", X"FE", X"FE"), (X"E9", X"E9", X"E9"), (X"BC", X"BC", X"BC"), (X"88", X"88", X"88"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"9E", X"9E", X"9E"), (X"9E", X"9E", X"9E"), (X"9E", X"9E", X"9E"), (X"9E", X"9E", X"9E"), (X"9E", X"9E", X"9E"), (X"9E", X"9E", X"9E"), (X"C5", X"C5", X"C5"), (X"DF", X"DC", X"DD"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"DE", X"DC", X"DC"), (X"D5", X"DC", X"D9"), (X"B9", X"C3", X"BF"), (X"B9", X"C3", X"BF"), (X"B9", X"C3", X"BF"), (X"B9", X"C3", X"BF"), (X"B9", X"C3", X"BF"), (X"B9", X"C3", X"BF"), (X"B9", X"C3", X"BF"), (X"B9", X"C3", X"BF"), (X"B9", X"C3", X"BF"), (X"D3", X"DD", X"DA"), (X"CD", X"D1", X"DA"), (X"BC", X"BF", X"C9"), (X"BC", X"BF", X"C9"), (X"BC", X"BF", X"C9"), (X"BC", X"BF", X"C9"), (X"BC", X"BF", X"C9"), (X"BC", X"BF", X"C9"), (X"BC", X"BF", X"C9"), (X"BC", X"BF", X"C9"), (X"BC", X"BF", X"C9"), (X"E3", X"E4", X"E8"), (X"D1", X"D1", X"D1"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"E8", X"E8", X"E8"), (X"CE", X"CE", X"CE"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"EB", X"EB", X"EB"), (X"CA", X"CA", X"CA"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"EE", X"EE", X"EE"), (X"D4", X"D4", X"D4"), (X"D6", X"D6", X"D6"), (X"F9", X"F9", X"F9"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B1", X"B1", X"B1"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"A3", X"A3", X"A3"), (X"AB", X"AB", X"AB"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FA", X"FA", X"FA"), (X"D8", X"D8", X"D8"), (X"D2", X"D2", X"D2"), (X"F1", X"F1", X"F1"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"C7", X"C7", X"C7"), (X"EE", X"EE", X"EE"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"CA", X"CA", X"CA"), (X"EB", X"EB", X"EB"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"CD", X"CD", X"CD"), (X"E7", X"E8", X"EC"), (X"BC", X"BF", X"C9"), (X"BC", X"BF", X"C9"), (X"BC", X"BF", X"C9"), (X"BC", X"BF", X"C9"), (X"BC", X"BF", X"C9"), (X"BC", X"BF", X"C9"), (X"BC", X"BF", X"C9"), (X"BC", X"BF", X"C9"), (X"BC", X"BF", X"C9"), (X"CA", X"CE", X"D7"), (X"DC", X"DF", X"D4"), (X"BF", X"C2", X"B4"), (X"BF", X"C2", X"B4"), (X"BF", X"C2", X"B4"), (X"BF", X"C2", X"B4"), (X"BF", X"C2", X"B4"), (X"BF", X"C2", X"B4"), (X"BF", X"C2", X"B4"), (X"BF", X"C2", X"B4"), (X"BF", X"C2", X"B4"), (X"D5", X"D7", X"CE"), (X"E0", X"E0", X"E3"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"D9", X"D8", X"DC"), (X"CB", X"CB", X"CB"), (X"9E", X"9E", X"9E"), (X"9E", X"9E", X"9E"), (X"9E", X"9E", X"9E"), (X"9E", X"9E", X"9E"), (X"9E", X"9E", X"9E"), (X"9E", X"9E", X"9E"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7C", X"7C", X"7C"), (X"A0", X"A0", X"A0"), (X"F1", X"F1", X"F1"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"26", X"26", X"26"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"16", X"16", X"16"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F5", X"F5", X"F5"), (X"A4", X"A4", X"A4"), (X"7C", X"7C", X"7C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"9F", X"9F", X"9F"), (X"E2", X"E2", X"E2"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"26", X"26", X"26"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"16", X"16", X"16"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"E6", X"E6", X"E6"), (X"A3", X"A3", X"A3"), (X"7B", X"7B", X"7B"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"94", X"94", X"94"), (X"DD", X"DD", X"DD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"26", X"26", X"26"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"16", X"16", X"16"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"E1", X"E1", X"E1"), (X"98", X"98", X"98"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"C9", X"C9", X"C9"), (X"FE", X"FE", X"FE"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"26", X"26", X"26"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"16", X"16", X"16"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FE", X"FE", X"FE"), (X"CE", X"CE", X"CE"), (X"88", X"88", X"88"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7B", X"7B", X"7B"), (X"AA", X"AA", X"AA"), (X"F3", X"F3", X"F3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"26", X"26", X"26"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"16", X"16", X"16"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"7C", X"7C", X"7C"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"9F", X"9F", X"9F"), (X"D6", X"D6", X"D6"), (X"FE", X"FE", X"FE"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"26", X"26", X"26"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"16", X"16", X"16"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"DB", X"DB", X"DB"), (X"9D", X"9D", X"9D"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DA", X"DA", X"DA"), (X"F9", X"F9", X"F9"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"26", X"26", X"26"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"16", X"16", X"16"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F9", X"F9", X"F9"), (X"E2", X"E2", X"E2"), (X"7B", X"7B", X"7B"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7E", X"7E", X"7E"), (X"C4", X"C4", X"C4"), (X"FE", X"FE", X"FE"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"26", X"26", X"26"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"16", X"16", X"16"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FE", X"FE", X"FE"), (X"CA", X"CA", X"CA"), (X"80", X"80", X"80"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B8", X"B8", X"B8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B7", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"88", X"88", X"88"), (X"DF", X"DF", X"DF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"26", X"26", X"26"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"16", X"16", X"16"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"E4", X"E4", X"E4"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C0"), (X"7A", X"7A", X"7B"), (X"7A", X"7A", X"7B"), (X"7A", X"7A", X"7B"), (X"7A", X"7A", X"7B"), (X"7A", X"7A", X"7B"), (X"7A", X"7A", X"7B"), (X"7A", X"7A", X"7B"), (X"7A", X"7A", X"7B"), (X"7A", X"7A", X"7B"), (X"B0", X"B0", X"B0"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"96", X"96", X"96"), (X"F0", X"F0", X"F0"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"26", X"26", X"26"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"16", X"16", X"16"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F4", X"F4", X"F4"), (X"9B", X"9B", X"9B"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"D6", X"D6", X"D6"), (X"D6", X"D6", X"D6"), (X"D6", X"D6", X"D6"), (X"D6", X"D6", X"D6"), (X"D6", X"D6", X"D6"), (X"D6", X"D6", X"D6"), (X"E6", X"E6", X"E6"), (X"DC", X"DE", X"DD"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"DB", X"DD", X"DC"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"D1", X"D1", X"D1"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"E8", X"E8", X"E8"), (X"CE", X"CE", X"CE"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"8E", X"8E", X"8E"), (X"8D", X"8D", X"8D"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"E9", X"E9", X"E9"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B0", X"B0", X"B0"), (X"F1", X"F1", X"F1"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"81", X"81", X"81"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"78", X"78", X"78"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"EF", X"EF", X"EF"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"90", X"90", X"90"), (X"8A", X"8A", X"8A"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"CA", X"CA", X"CA"), (X"EB", X"EB", X"EB"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"CD", X"CD", X"CD"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"E0", X"E1", X"DE"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"D9", X"DA", X"D6"), (X"E9", X"E9", X"E9"), (X"D6", X"D6", X"D6"), (X"D6", X"D6", X"D6"), (X"D6", X"D6", X"D6"), (X"D6", X"D6", X"D6"), (X"D6", X"D6", X"D6"), (X"D6", X"D6", X"D6"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"4A", X"4A", X"4A"), (X"03", X"03", X"03"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"CA", X"CA", X"CA"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"44", X"44", X"44"), (X"DD", X"DD", X"DD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"DA", X"DA", X"DA"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"02", X"02"), (X"43", X"43", X"43"), (X"79", X"79", X"79"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"79", X"79", X"79"), (X"44", X"44", X"44"), (X"02", X"02", X"02"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"CA", X"CA", X"CA"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"44", X"44", X"44"), (X"DD", X"DD", X"DD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"DA", X"DA", X"DA"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"01", X"01", X"01"), (X"3D", X"3D", X"3D"), (X"79", X"79", X"79"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"42", X"42", X"42"), (X"01", X"01", X"01"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"CA", X"CA", X"CA"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"44", X"44", X"44"), (X"DD", X"DD", X"DD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"DA", X"DA", X"DA"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"01", X"01", X"01"), (X"3B", X"3B", X"3B"), (X"79", X"79", X"79"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"45", X"45", X"45"), (X"01", X"01", X"01"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"CA", X"CA", X"CA"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"44", X"44", X"44"), (X"DD", X"DD", X"DD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"DA", X"DA", X"DA"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"01", X"01", X"01"), (X"3D", X"3D", X"3D"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"68", X"68", X"68"), (X"02", X"02", X"02"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"CA", X"CA", X"CA"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"44", X"44", X"44"), (X"DD", X"DD", X"DD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"DA", X"DA", X"DA"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"01", X"01", X"01"), (X"59", X"59", X"59"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"06", X"06", X"06"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"CA", X"CA", X"CA"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"44", X"44", X"44"), (X"DD", X"DD", X"DD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"DA", X"DA", X"DA"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"02", X"02"), (X"82", X"82", X"82"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"63", X"63", X"63"), (X"08", X"08", X"08"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"CA", X"CA", X"CA"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"44", X"44", X"44"), (X"DD", X"DD", X"DD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"DA", X"DA", X"DA"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"06", X"06", X"06"), (X"5D", X"5D", X"5D"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"6F", X"6F", X"6F"), (X"10", X"10", X"10"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"CA", X"CA", X"CA"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"44", X"44", X"44"), (X"DD", X"DD", X"DD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"DA", X"DA", X"DA"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"0D", X"0D", X"0D"), (X"6B", X"6B", X"6B"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"77", X"77", X"77"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"CA", X"CA", X"CA"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"44", X"44", X"44"), (X"DD", X"DD", X"DD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"DA", X"DA", X"DA"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"1C", X"1C", X"1C"), (X"75", X"75", X"75"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3E", X"97", X"82"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"B8", X"C7", X"EE"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"3C", X"3C", X"3C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"CA", X"CA", X"CA"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"44", X"44", X"44"), (X"DD", X"DD", X"DD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"DA", X"DA", X"DA"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"34", X"34", X"34"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"C3", X"CF", X"F0"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"57", X"7A", X"D6"), (X"75", X"8D", X"29"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"C5", X"C5", X"C5"), (X"C5", X"C5", X"C5"), (X"C5", X"C5", X"C5"), (X"C5", X"C5", X"C5"), (X"C5", X"C5", X"C5"), (X"C5", X"C5", X"C5"), (X"DC", X"DC", X"DC"), (X"DC", X"DD", X"DD"), (X"BE", X"C0", X"BF"), (X"BE", X"C0", X"BF"), (X"BE", X"C0", X"BF"), (X"BE", X"C0", X"BF"), (X"BE", X"C0", X"BF"), (X"BE", X"C0", X"BF"), (X"BE", X"C0", X"BF"), (X"BE", X"C0", X"BF"), (X"BE", X"C0", X"BF"), (X"DC", X"DD", X"DC"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"8B", X"C2", X"B1"), (X"C3", X"CB", X"E0"), (X"B7", X"BF", X"D4"), (X"B7", X"BF", X"D4"), (X"B7", X"BF", X"D4"), (X"B7", X"BF", X"D4"), (X"B7", X"BF", X"D4"), (X"B7", X"BF", X"D4"), (X"B7", X"BF", X"D4"), (X"B7", X"BF", X"D4"), (X"B7", X"BF", X"D4"), (X"E1", X"E4", X"ED"), (X"D1", X"D1", X"D1"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"B6", X"B6", X"B6"), (X"64", X"64", X"64"), (X"62", X"62", X"62"), (X"62", X"62", X"62"), (X"62", X"62", X"62"), (X"62", X"62", X"62"), (X"62", X"62", X"62"), (X"55", X"55", X"55"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2B", X"2B", X"2B"), (X"62", X"62", X"62"), (X"62", X"62", X"62"), (X"62", X"62", X"62"), (X"62", X"62", X"62"), (X"62", X"62", X"62"), (X"C4", X"C4", X"C4"), (X"DE", X"DE", X"DE"), (X"96", X"96", X"96"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"21", X"21", X"21"), (X"6C", X"6C", X"6C"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"86", X"86", X"86"), (X"DA", X"DA", X"DA"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"BC", X"BC", X"BC"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"BD", X"BD", X"BD"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"80", X"80", X"80"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"97", X"97", X"97"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"A6", X"A6", X"A6"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"7D", X"7D", X"7D"), (X"7F", X"7F", X"7F"), (X"D1", X"D1", X"D1"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"DE", X"DE", X"DE"), (X"CB", X"CB", X"CB"), (X"7D", X"7D", X"7D"), (X"6B", X"6B", X"6B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"30", X"30", X"30"), (X"62", X"62", X"62"), (X"62", X"62", X"62"), (X"62", X"62", X"62"), (X"62", X"62", X"62"), (X"62", X"62", X"62"), (X"62", X"62", X"62"), (X"62", X"62", X"62"), (X"14", X"14", X"14"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"01", X"01", X"01"), (X"7F", X"7F", X"7F"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"CD", X"CD", X"CD"), (X"E5", X"E8", X"F0"), (X"B7", X"BF", X"D4"), (X"B7", X"BF", X"D4"), (X"B7", X"BF", X"D4"), (X"B7", X"BF", X"D4"), (X"B7", X"BF", X"D4"), (X"B7", X"BF", X"D4"), (X"B7", X"BF", X"D4"), (X"B7", X"BF", X"D4"), (X"B7", X"BF", X"D4"), (X"C1", X"C9", X"DE"), (X"B5", X"C1", X"7F"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"E0", X"E1", X"DF"), (X"BF", X"C0", X"BD"), (X"BF", X"C0", X"BD"), (X"BF", X"C0", X"BD"), (X"BF", X"C0", X"BD"), (X"BF", X"C0", X"BD"), (X"BF", X"C0", X"BD"), (X"BF", X"C0", X"BD"), (X"BF", X"C0", X"BD"), (X"BF", X"C0", X"BD"), (X"D9", X"DA", X"D8"), (X"E0", X"E0", X"E0"), (X"C5", X"C5", X"C5"), (X"C5", X"C5", X"C5"), (X"C5", X"C5", X"C5"), (X"C5", X"C5", X"C5"), (X"C5", X"C5", X"C5"), (X"C5", X"C5", X"C5"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"6F", X"6F", X"6F"), (X"A5", X"A5", X"A5"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"A6", X"A6", X"A6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"54", X"54", X"54"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"32", X"32", X"32"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"11", X"11", X"11"), (X"B7", X"B7", X"B7"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"7C", X"7C", X"7C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"7F", X"7F", X"7F"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"06", X"06", X"06"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"33", X"33", X"33"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"51", X"51", X"51"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"A5", X"A5", X"A5"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"9A", X"9A", X"9A"), (X"01", X"01", X"01"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"5D", X"5D", X"5D"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"27", X"27", X"27"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"15", X"15", X"15"), (X"82", X"82", X"82"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"2B", X"2B", X"2B"), (X"9E", X"9E", X"9E"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"A6", X"A6", X"A6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"54", X"54", X"54"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"32", X"32", X"32"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"11", X"11", X"11"), (X"B7", X"B7", X"B7"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"7C", X"7C", X"7C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"7F", X"7F", X"7F"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"06", X"06", X"06"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"33", X"33", X"33"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"51", X"51", X"51"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"A5", X"A5", X"A5"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"9A", X"9A", X"9A"), (X"01", X"01", X"01"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"5D", X"5D", X"5D"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"27", X"27", X"27"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"14", X"14", X"14"), (X"AB", X"AB", X"AB"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"54", X"54", X"54"), (X"01", X"01", X"01"), (X"9E", X"9E", X"9E"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"A6", X"A6", X"A6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"54", X"54", X"54"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"32", X"32", X"32"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"11", X"11", X"11"), (X"B7", X"B7", X"B7"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"7C", X"7C", X"7C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"7F", X"7F", X"7F"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"06", X"06", X"06"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"33", X"33", X"33"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"51", X"51", X"51"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"A5", X"A5", X"A5"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"9A", X"9A", X"9A"), (X"01", X"01", X"01"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"5D", X"5D", X"5D"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"27", X"27", X"27"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"14", X"14", X"14"), (X"BF", X"BF", X"BF"), (X"93", X"93", X"93"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"74", X"74", X"74"), (X"0F", X"0F", X"0F"), (X"00", X"00", X"00"), (X"9E", X"9E", X"9E"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"A6", X"A6", X"A6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"54", X"54", X"54"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"32", X"32", X"32"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"11", X"11", X"11"), (X"B7", X"B7", X"B7"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"7C", X"7C", X"7C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"7F", X"7F", X"7F"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"06", X"06", X"06"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"33", X"33", X"33"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"51", X"51", X"51"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"A5", X"A5", X"A5"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"9A", X"9A", X"9A"), (X"01", X"01", X"01"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"5D", X"5D", X"5D"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"27", X"27", X"27"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"14", X"14", X"14"), (X"BF", X"BF", X"BF"), (X"B9", X"B9", X"B9"), (X"80", X"80", X"80"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"3A", X"3A", X"3A"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"9E", X"9E", X"9E"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"A6", X"A6", X"A6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"54", X"54", X"54"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"32", X"32", X"32"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"11", X"11", X"11"), (X"B7", X"B7", X"B7"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"7C", X"7C", X"7C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"7F", X"7F", X"7F"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"06", X"06", X"06"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"33", X"33", X"33"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"51", X"51", X"51"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"A5", X"A5", X"A5"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"9A", X"9A", X"9A"), (X"01", X"01", X"01"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"5D", X"5D", X"5D"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"27", X"27", X"27"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"14", X"14", X"14"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"A2", X"A2", X"A2"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"6A", X"6A", X"6A"), (X"04", X"04", X"04"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"9E", X"9E", X"9E"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"A6", X"A6", X"A6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"54", X"54", X"54"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"32", X"32", X"32"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"11", X"11", X"11"), (X"B7", X"B7", X"B7"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"7C", X"7C", X"7C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"7F", X"7F", X"7F"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"06", X"06", X"06"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"33", X"33", X"33"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"51", X"51", X"51"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"A5", X"A5", X"A5"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"9A", X"9A", X"9A"), (X"01", X"01", X"01"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"5D", X"5D", X"5D"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"27", X"27", X"27"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"14", X"14", X"14"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BD", X"BD", X"BD"), (X"87", X"87", X"87"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"79", X"79", X"79"), (X"29", X"29", X"29"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"9E", X"9E", X"9E"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"A6", X"A6", X"A6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"54", X"54", X"54"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"32", X"32", X"32"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"11", X"11", X"11"), (X"B7", X"B7", X"B7"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"7C", X"7C", X"7C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"7F", X"7F", X"7F"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"06", X"06", X"06"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"33", X"33", X"33"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"51", X"51", X"51"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"A5", X"A5", X"A5"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"9A", X"9A", X"9A"), (X"01", X"01", X"01"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"5D", X"5D", X"5D"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"27", X"27", X"27"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"14", X"14", X"14"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"AB", X"AB", X"AB"), (X"7B", X"7B", X"7B"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"60", X"60", X"60"), (X"02", X"02", X"02"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"9E", X"9E", X"9E"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"A6", X"A6", X"A6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"54", X"54", X"54"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"32", X"32", X"32"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"11", X"11", X"11"), (X"B7", X"B7", X"B7"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"7C", X"7C", X"7C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"7F", X"7F", X"7F"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"06", X"06", X"06"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"33", X"33", X"33"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"51", X"51", X"51"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"A5", X"A5", X"A5"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"9A", X"9A", X"9A"), (X"01", X"01", X"01"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"5D", X"5D", X"5D"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"27", X"27", X"27"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"14", X"14", X"14"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BE", X"BE", X"BE"), (X"8C", X"8C", X"8C"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"24", X"24", X"24"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"9E", X"9E", X"9E"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"A6", X"A6", X"A6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"54", X"54", X"54"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"32", X"32", X"32"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"11", X"11", X"11"), (X"B7", X"B7", X"B7"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"7C", X"7C", X"7C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"7F", X"7F", X"7F"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"06", X"06", X"06"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"33", X"33", X"33"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"51", X"51", X"51"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"A5", X"A5", X"A5"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"9A", X"9A", X"9A"), (X"01", X"01", X"01"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"5D", X"5D", X"5D"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"27", X"27", X"27"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"14", X"14", X"14"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"AE", X"AE", X"AE"), (X"99", X"99", X"99"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"87", X"87", X"87"), (X"02", X"02", X"02"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"9E", X"9E", X"9E"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"A6", X"A6", X"A6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"54", X"54", X"54"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"32", X"32", X"32"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"11", X"11", X"11"), (X"B7", X"B7", X"B7"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"7C", X"7C", X"7C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"7F", X"7F", X"7F"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"06", X"06", X"06"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"33", X"33", X"33"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"51", X"51", X"51"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"A5", X"A5", X"A5"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"9A", X"9A", X"9A"), (X"01", X"01", X"01"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"5D", X"5D", X"5D"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"27", X"27", X"27"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"14", X"14", X"14"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BE", X"BE", X"BE"), (X"AA", X"AA", X"AA"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"B0", X"B0", X"B0"), (X"B0", X"B0", X"B0"), (X"B0", X"B0", X"B0"), (X"B0", X"B0", X"B0"), (X"B0", X"B0", X"B0"), (X"B0", X"B0", X"B0"), (X"D0", X"D0", X"D0"), (X"DF", X"DC", X"DD"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"DE", X"DC", X"DC"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"D5", X"D5", X"D5"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"E4", X"E4", X"E4"), (X"A3", X"A3", X"50"), (X"6D", X"6D", X"00"), (X"6D", X"6D", X"00"), (X"6D", X"6D", X"00"), (X"6D", X"6D", X"00"), (X"6D", X"6D", X"00"), (X"B1", X"B1", X"44"), (X"BF", X"BF", X"52"), (X"BF", X"BF", X"52"), (X"BF", X"BF", X"52"), (X"BF", X"BF", X"52"), (X"BF", X"BF", X"52"), (X"BF", X"BF", X"52"), (X"B4", X"B4", X"47"), (X"6D", X"6D", X"00"), (X"6D", X"6D", X"00"), (X"1D", X"6D", X"50"), (X"00", X"6D", X"6D"), (X"00", X"6D", X"6D"), (X"00", X"6D", X"6D"), (X"00", X"6D", X"6D"), (X"24", X"91", X"91"), (X"52", X"BF", X"BF"), (X"52", X"BF", X"BF"), (X"52", X"BF", X"BF"), (X"52", X"BF", X"BF"), (X"52", X"BF", X"BF"), (X"52", X"BF", X"BF"), (X"52", X"BF", X"BF"), (X"15", X"82", X"82"), (X"00", X"6D", X"6D"), (X"00", X"6D", X"6D"), (X"00", X"6D", X"6D"), (X"00", X"6D", X"6D"), (X"00", X"6D", X"6D"), (X"00", X"6D", X"6D"), (X"08", X"75", X"75"), (X"4E", X"BB", X"BB"), (X"52", X"BF", X"62"), (X"52", X"BF", X"52"), (X"52", X"BF", X"52"), (X"52", X"BF", X"52"), (X"52", X"BF", X"52"), (X"52", X"BF", X"52"), (X"35", X"A2", X"35"), (X"00", X"6D", X"00"), (X"00", X"6D", X"00"), (X"00", X"6D", X"00"), (X"00", X"6D", X"00"), (X"00", X"6D", X"00"), (X"00", X"6D", X"00"), (X"00", X"6D", X"00"), (X"36", X"A3", X"36"), (X"52", X"BF", X"52"), (X"52", X"BF", X"52"), (X"52", X"BF", X"52"), (X"52", X"BF", X"52"), (X"52", X"BF", X"52"), (X"52", X"BF", X"52"), (X"52", X"BF", X"52"), (X"6C", X"06", X"6C"), (X"6D", X"00", X"6D"), (X"6D", X"00", X"6D"), (X"6D", X"00", X"6D"), (X"6D", X"00", X"6D"), (X"6D", X"00", X"6D"), (X"6D", X"00", X"6D"), (X"83", X"16", X"83"), (X"BF", X"52", X"BF"), (X"BF", X"52", X"BF"), (X"BF", X"52", X"BF"), (X"BF", X"52", X"BF"), (X"BF", X"52", X"BF"), (X"BF", X"52", X"BF"), (X"BF", X"52", X"BF"), (X"90", X"23", X"90"), (X"6D", X"00", X"6D"), (X"6D", X"00", X"6D"), (X"6D", X"00", X"6D"), (X"6D", X"00", X"6D"), (X"6D", X"00", X"6D"), (X"6D", X"00", X"64"), (X"6E", X"01", X"01"), (X"B4", X"47", X"47"), (X"BF", X"52", X"52"), (X"BF", X"52", X"52"), (X"BF", X"52", X"52"), (X"BF", X"52", X"52"), (X"BF", X"52", X"52"), (X"BF", X"52", X"52"), (X"AF", X"42", X"42"), (X"6D", X"00", X"00"), (X"6D", X"00", X"00"), (X"6D", X"00", X"00"), (X"6D", X"00", X"00"), (X"6D", X"00", X"00"), (X"6D", X"00", X"00"), (X"6D", X"00", X"00"), (X"95", X"28", X"28"), (X"BF", X"52", X"52"), (X"BF", X"52", X"52"), (X"BF", X"52", X"52"), (X"BF", X"52", X"52"), (X"A9", X"52", X"68"), (X"52", X"52", X"BF"), (X"52", X"52", X"BF"), (X"11", X"11", X"7E"), (X"00", X"00", X"6D"), (X"00", X"00", X"6D"), (X"00", X"00", X"6D"), (X"00", X"00", X"6D"), (X"00", X"00", X"6D"), (X"00", X"00", X"6D"), (X"08", X"08", X"75"), (X"52", X"52", X"BF"), (X"52", X"52", X"BF"), (X"52", X"52", X"BF"), (X"52", X"52", X"BF"), (X"52", X"52", X"BF"), (X"70", X"70", X"CA"), (X"E7", X"E7", X"E8"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"D1", X"D1", X"D1"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"E0", X"E0", X"E3"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"D9", X"D8", X"DC"), (X"D5", X"D5", X"D5"), (X"B0", X"B0", X"B0"), (X"B0", X"B0", X"B0"), (X"B0", X"B0", X"B0"), (X"B0", X"B0", X"B0"), (X"B0", X"B0", X"B0"), (X"B0", X"B0", X"B0"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BE", X"BE", X"A3"), (X"C1", X"C1", X"08"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"B9", X"06", X"B9"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"04", X"04", X"C0"), (X"A0", X"A0", X"C3"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"78", X"7B", X"7A"), (X"78", X"7B", X"7A"), (X"78", X"7B", X"7A"), (X"78", X"7B", X"7A"), (X"78", X"7B", X"7A"), (X"78", X"7B", X"7A"), (X"78", X"7B", X"7A"), (X"78", X"7B", X"7A"), (X"78", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"AB", X"AB", X"45"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"B9", X"06", X"B9"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"3D", X"3D", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BE"), (X"7A", X"7B", X"77"), (X"7A", X"7B", X"77"), (X"7A", X"7B", X"77"), (X"7A", X"7B", X"77"), (X"7A", X"7B", X"77"), (X"7A", X"7B", X"77"), (X"7A", X"7B", X"77"), (X"7A", X"7B", X"77"), (X"7A", X"7B", X"77"), (X"B0", X"B0", X"AE"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7D", X"7D", X"75"), (X"B8", X"B8", X"0C"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"B9", X"06", X"B9"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"06", X"06", X"BB"), (X"73", X"73", X"7E"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"91", X"91", X"51"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"B9", X"06", X"B9"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"49", X"49", X"96"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"AA", X"AA", X"24"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"B9", X"06", X"B9"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"1D", X"1D", X"AE"), (X"79", X"79", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"80", X"80", X"6F"), (X"BD", X"BD", X"04"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"B9", X"06", X"B9"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"01", X"01", X"BE"), (X"6A", X"6A", X"83"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"95", X"95", X"4A"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"B9", X"06", X"B9"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"43", X"43", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"AB", X"AB", X"23"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"B9", X"06", X"B9"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"1C", X"1C", X"AF"), (X"79", X"79", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7D", X"7D", X"74"), (X"BC", X"BC", X"04"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"B9", X"06", X"B9"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"03", X"03", X"BD"), (X"6E", X"6E", X"81"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8E", X"8E", X"56"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"B9", X"06", X"B9"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"4F", X"4F", X"92"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"E3", X"E3", X"E3"), (X"E3", X"E3", X"E3"), (X"E3", X"E3", X"E3"), (X"E3", X"E3", X"E3"), (X"E3", X"E3", X"E3"), (X"E3", X"E3", X"E3"), (X"EE", X"EE", X"EE"), (X"DC", X"DE", X"DD"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"DB", X"DD", X"DC"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"D5", X"D5", X"D5"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"C1", X"C1", X"57"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"B8", X"00"), (X"00", X"4E", X"00"), (X"00", X"47", X"00"), (X"00", X"47", X"00"), (X"00", X"47", X"00"), (X"41", X"88", X"41"), (X"8F", X"4D", X"8F"), (X"47", X"00", X"47"), (X"47", X"00", X"47"), (X"47", X"00", X"47"), (X"49", X"00", X"49"), (X"B5", X"00", X"B5"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"4B", X"4B", X"C1"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"D1", X"D1", X"D1"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"E0", X"E1", X"DE"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"D9", X"DA", X"D6"), (X"F0", X"F0", X"F0"), (X"E3", X"E3", X"E3"), (X"E3", X"E3", X"E3"), (X"E3", X"E3", X"E3"), (X"E3", X"E3", X"E3"), (X"E3", X"E3", X"E3"), (X"E3", X"E3", X"E3"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7B", X"7B", X"79"), (X"B1", X"B1", X"19"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"B4", X"00"), (X"00", X"0A", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"00", X"02"), (X"B0", X"00", X"B0"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"12", X"12", X"B5"), (X"78", X"78", X"7B"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7E", X"7E", X"72"), (X"BD", X"BD", X"04"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"B4", X"00"), (X"00", X"0A", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"00", X"02"), (X"B0", X"00", X"B0"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"02", X"02", X"BE"), (X"6C", X"6C", X"82"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B8", X"B8", X"B8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B7", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"5B"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"B4", X"00"), (X"00", X"0A", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"00", X"02"), (X"B0", X"00", X"B0"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"54", X"54", X"8F"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"C0", X"BF"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"B0", X"B0", X"AF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"99", X"99", X"43"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"B4", X"00"), (X"00", X"0A", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"00", X"02"), (X"B0", X"00", X"B0"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"3B", X"3B", X"9D"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A5", X"A5", X"2D"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"B4", X"00"), (X"00", X"0A", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"00", X"02"), (X"B0", X"00", X"B0"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"25", X"25", X"AA"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B1", X"B1", X"19"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"B4", X"00"), (X"00", X"0A", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"00", X"02"), (X"B0", X"00", X"B0"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"11", X"11", X"B5"), (X"79", X"79", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7D", X"7D", X"75"), (X"B9", X"B9", X"0B"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"B4", X"00"), (X"00", X"0A", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"00", X"02"), (X"B0", X"00", X"B0"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"07", X"07", X"BB"), (X"71", X"71", X"7F"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"81", X"81", X"6E"), (X"BE", X"BE", X"02"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"B4", X"00"), (X"00", X"0A", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"00", X"02"), (X"B0", X"00", X"B0"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"01", X"01", X"BE"), (X"67", X"67", X"85"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"88", X"88", X"61"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"B4", X"00"), (X"00", X"0A", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"00", X"02"), (X"B0", X"00", X"B0"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"59", X"59", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8F", X"8F", X"54"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"33", X"BF", X"8C"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"BF"), (X"00", X"BF", X"1D"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"BF", X"00"), (X"00", X"B4", X"00"), (X"00", X"0A", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"00", X"02"), (X"B0", X"00", X"B0"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"BF"), (X"BF", X"00", X"AE"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"98", X"00", X"27"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"00", X"00", X"BF"), (X"4C", X"4C", X"94"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"92", X"92", X"92"), (X"92", X"92", X"92"), (X"92", X"92", X"92"), (X"92", X"92", X"92"), (X"92", X"92", X"92"), (X"92", X"92", X"92"), (X"BE", X"BE", X"BE"), (X"DF", X"DC", X"DD"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"C2", X"BE", X"BF"), (X"DE", X"DC", X"DC"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"D5", X"D5", X"D5"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"8A", X"8A", X"74"), (X"3B", X"3B", X"00"), (X"3B", X"3B", X"00"), (X"3B", X"3B", X"00"), (X"3B", X"3B", X"00"), (X"A1", X"A1", X"66"), (X"6E", X"6E", X"33"), (X"3B", X"3B", X"00"), (X"3B", X"3B", X"00"), (X"3B", X"3B", X"00"), (X"3B", X"3B", X"00"), (X"3B", X"3B", X"00"), (X"3B", X"3B", X"00"), (X"3B", X"3B", X"00"), (X"3B", X"3B", X"00"), (X"3B", X"3B", X"00"), (X"AB", X"AB", X"70"), (X"64", X"64", X"29"), (X"3B", X"3B", X"00"), (X"3B", X"3B", X"00"), (X"3B", X"3B", X"00"), (X"3B", X"3B", X"00"), (X"10", X"3B", X"2B"), (X"00", X"3B", X"3B"), (X"00", X"3B", X"3B"), (X"00", X"3B", X"3B"), (X"00", X"3B", X"3B"), (X"7A", X"B6", X"B6"), (X"1E", X"5A", X"5A"), (X"00", X"3B", X"3B"), (X"00", X"3B", X"3B"), (X"00", X"3B", X"3B"), (X"00", X"3B", X"3B"), (X"00", X"3B", X"3B"), (X"00", X"3B", X"3B"), (X"00", X"3B", X"3B"), (X"00", X"3B", X"3B"), (X"00", X"3B", X"3B"), (X"81", X"BD", X"BD"), (X"17", X"53", X"53"), (X"00", X"3B", X"3B"), (X"00", X"3B", X"3B"), (X"00", X"3B", X"3B"), (X"00", X"3B", X"3B"), (X"00", X"3B", X"09"), (X"00", X"3B", X"00"), (X"00", X"3B", X"00"), (X"00", X"3B", X"00"), (X"00", X"3B", X"00"), (X"88", X"C4", X"88"), (X"10", X"4C", X"10"), (X"00", X"3B", X"00"), (X"00", X"3B", X"00"), (X"00", X"3B", X"00"), (X"00", X"3B", X"00"), (X"00", X"3B", X"00"), (X"00", X"3B", X"00"), (X"00", X"3B", X"00"), (X"00", X"3B", X"00"), (X"00", X"3B", X"00"), (X"8F", X"C7", X"8F"), (X"0A", X"0D", X"0A"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"02", X"03"), (X"CA", X"94", X"CA"), (X"3E", X"03", X"3E"), (X"3B", X"00", X"3B"), (X"3B", X"00", X"3B"), (X"3B", X"00", X"3B"), (X"3B", X"00", X"3B"), (X"3B", X"00", X"3B"), (X"3B", X"00", X"3B"), (X"3B", X"00", X"3B"), (X"3B", X"00", X"3B"), (X"44", X"09", X"44"), (X"CB", X"8F", X"CB"), (X"3B", X"00", X"3B"), (X"3B", X"00", X"3B"), (X"3B", X"00", X"3B"), (X"3B", X"00", X"3B"), (X"3B", X"00", X"36"), (X"3B", X"00", X"00"), (X"3B", X"00", X"00"), (X"3B", X"00", X"00"), (X"3B", X"00", X"00"), (X"4B", X"10", X"10"), (X"C4", X"89", X"89"), (X"3B", X"00", X"00"), (X"3B", X"00", X"00"), (X"3B", X"00", X"00"), (X"3B", X"00", X"00"), (X"3B", X"00", X"00"), (X"3B", X"00", X"00"), (X"3B", X"00", X"00"), (X"3B", X"00", X"00"), (X"3B", X"00", X"00"), (X"52", X"17", X"17"), (X"BD", X"82", X"82"), (X"3B", X"00", X"00"), (X"3B", X"00", X"00"), (X"3B", X"00", X"00"), (X"3B", X"00", X"00"), (X"2F", X"00", X"0C"), (X"00", X"00", X"3B"), (X"00", X"00", X"3B"), (X"00", X"00", X"3B"), (X"00", X"00", X"3B"), (X"1E", X"1E", X"59"), (X"7B", X"7B", X"B6"), (X"00", X"00", X"3B"), (X"00", X"00", X"3B"), (X"00", X"00", X"3B"), (X"00", X"00", X"3B"), (X"00", X"00", X"3B"), (X"00", X"00", X"3B"), (X"00", X"00", X"3B"), (X"00", X"00", X"3B"), (X"00", X"00", X"3B"), (X"28", X"28", X"63"), (X"71", X"71", X"AC"), (X"00", X"00", X"3B"), (X"00", X"00", X"3B"), (X"00", X"00", X"3B"), (X"00", X"00", X"3B"), (X"68", X"68", X"81"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"D1", X"D1", X"D1"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"E0", X"E0", X"E3"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"BF", X"BE", X"C4"), (X"D9", X"D8", X"DC"), (X"C5", X"C5", X"C5"), (X"92", X"92", X"92"), (X"92", X"92", X"92"), (X"92", X"92", X"92"), (X"92", X"92", X"92"), (X"92", X"92", X"92"), (X"92", X"92", X"92"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"40", X"40", X"40"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"93", X"93", X"93"), (X"4A", X"4A", X"4A"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"A2", X"A2", X"A2"), (X"3B", X"3B", X"3B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"B1", X"B1", X"B1"), (X"2C", X"2C", X"2C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"C5", X"C5", X"C5"), (X"18", X"18", X"18"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"D0", X"D0", X"D0"), (X"0E", X"0E", X"0E"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"D6", X"D6", X"D6"), (X"04", X"04", X"04"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"0D", X"0D", X"0D"), (X"D0", X"D0", X"D0"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"17", X"17", X"17"), (X"C6", X"C6", X"C6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"21", X"21", X"21"), (X"BC", X"BC", X"BC"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2B", X"2B", X"2B"), (X"B2", X"B2", X"B2"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"3A", X"3A", X"3A"), (X"A3", X"A3", X"A3"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"39", X"39", X"39"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"39", X"39", X"39"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"93", X"93", X"93"), (X"4A", X"4A", X"4A"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"A2", X"A2", X"A2"), (X"3B", X"3B", X"3B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"B1", X"B1", X"B1"), (X"2C", X"2C", X"2C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"C5", X"C5", X"C5"), (X"18", X"18", X"18"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"D0", X"D0", X"D0"), (X"0E", X"0E", X"0E"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"D6", X"D6", X"D6"), (X"04", X"04", X"04"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"0D", X"0D", X"0D"), (X"D0", X"D0", X"D0"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"17", X"17", X"17"), (X"C6", X"C6", X"C6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"21", X"21", X"21"), (X"BC", X"BC", X"BC"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2B", X"2B", X"2B"), (X"B2", X"B2", X"B2"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"3A", X"3A", X"3A"), (X"A3", X"A3", X"A3"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"32", X"32", X"32"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"34", X"34", X"34"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"93", X"93", X"93"), (X"4A", X"4A", X"4A"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"A2", X"A2", X"A2"), (X"3B", X"3B", X"3B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"B1", X"B1", X"B1"), (X"2C", X"2C", X"2C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"C5", X"C5", X"C5"), (X"18", X"18", X"18"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"D0", X"D0", X"D0"), (X"0E", X"0E", X"0E"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"D6", X"D6", X"D6"), (X"04", X"04", X"04"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"0D", X"0D", X"0D"), (X"D0", X"D0", X"D0"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"17", X"17", X"17"), (X"C6", X"C6", X"C6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"21", X"21", X"21"), (X"BC", X"BC", X"BC"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2B", X"2B", X"2B"), (X"B2", X"B2", X"B2"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"3A", X"3A", X"3A"), (X"A3", X"A3", X"A3"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2C", X"2C", X"2C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"8C", X"C3", X"B0"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"3C", X"9A", X"7A"), (X"A1", X"CE", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"31", X"31", X"31"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"93", X"93", X"93"), (X"4A", X"4A", X"4A"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"A2", X"A2", X"A2"), (X"3B", X"3B", X"3B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"B1", X"B1", X"B1"), (X"2C", X"2C", X"2C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"C5", X"C5", X"C5"), (X"18", X"18", X"18"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"D0", X"D0", X"D0"), (X"0E", X"0E", X"0E"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"D6", X"D6", X"D6"), (X"04", X"04", X"04"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"0D", X"0D", X"0D"), (X"D0", X"D0", X"D0"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"17", X"17", X"17"), (X"C6", X"C6", X"C6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"21", X"21", X"21"), (X"BC", X"BC", X"BC"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2B", X"2B", X"2B"), (X"B2", X"B2", X"B2"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"3A", X"3A", X"3A"), (X"A3", X"A3", X"A3"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"29", X"29", X"29"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"D1", X"99"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"7A", X"90", X"0B"), (X"A8", X"B6", X"5F"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"A8", X"C0", X"B8"), (X"5C", X"89", X"7A"), (X"5C", X"89", X"7A"), (X"5C", X"89", X"7A"), (X"5C", X"89", X"7A"), (X"5C", X"89", X"7A"), (X"5C", X"89", X"7A"), (X"5C", X"89", X"7A"), (X"5C", X"89", X"7A"), (X"5C", X"89", X"7A"), (X"A7", X"BF", X"B7"), (X"9E", X"BA", X"B0"), (X"5B", X"8A", X"7A"), (X"5B", X"8A", X"7A"), (X"5B", X"8A", X"7A"), (X"5B", X"8A", X"7A"), (X"5B", X"8A", X"7A"), (X"5B", X"8A", X"7A"), (X"5B", X"8A", X"7A"), (X"5B", X"8A", X"7A"), (X"5B", X"8A", X"7A"), (X"B0", X"C7", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7F", X"7F", X"7F"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"CA", X"CA", X"CA"), (X"A6", X"A6", X"A6"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"D2", X"D2", X"D2"), (X"9F", X"9F", X"9F"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"D9", X"D9", X"D9"), (X"97", X"97", X"97"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"DE", X"DE", X"DE"), (X"93", X"93", X"93"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"E3", X"E3", X"E3"), (X"8E", X"8E", X"8E"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"E8", X"E8", X"E8"), (X"89", X"89", X"89"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"B4", X"B4", X"B4"), (X"BC", X"BC", X"BC"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"84", X"84", X"84"), (X"EB", X"EB", X"EB"), (X"84", X"84", X"84"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"89", X"89", X"89"), (X"E8", X"E8", X"E8"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"8D", X"8D", X"8D"), (X"E3", X"E3", X"E3"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"92", X"92", X"92"), (X"DE", X"DE", X"DE"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"97", X"97", X"97"), (X"D9", X"D9", X"D9"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"9E", X"9E", X"9E"), (X"D2", X"D2", X"D2"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"7F", X"7F", X"7F"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"CC", X"B0"), (X"7A", X"85", X"43"), (X"7A", X"85", X"43"), (X"7A", X"85", X"43"), (X"7A", X"85", X"43"), (X"7A", X"85", X"43"), (X"7A", X"85", X"43"), (X"7A", X"85", X"43"), (X"7A", X"85", X"43"), (X"7A", X"85", X"43"), (X"A8", X"AF", X"84"), (X"BF", X"C5", X"A6"), (X"7A", X"85", X"45"), (X"7A", X"85", X"45"), (X"7A", X"85", X"45"), (X"7A", X"85", X"45"), (X"7A", X"85", X"45"), (X"7A", X"85", X"45"), (X"7A", X"85", X"45"), (X"7A", X"85", X"45"), (X"7A", X"85", X"45"), (X"B0", X"B6", X"90"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"31", X"31", X"31"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"94", X"94", X"94"), (X"4C", X"4C", X"4C"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"A3", X"A3", X"A3"), (X"3D", X"3D", X"3D"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"B2", X"B2", X"B2"), (X"2E", X"2E", X"2E"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"BC", X"BC", X"BC"), (X"24", X"24", X"24"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"C6", X"C6", X"C6"), (X"1A", X"1A", X"1A"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"D0", X"D0", X"D0"), (X"10", X"10", X"10"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"68", X"68", X"68"), (X"78", X"78", X"78"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"05", X"05", X"05"), (X"D7", X"D7", X"D7"), (X"06", X"06", X"06"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"0F", X"0F", X"0F"), (X"D1", X"D1", X"D1"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"19", X"19", X"19"), (X"C7", X"C7", X"C7"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"23", X"23", X"23"), (X"BD", X"BD", X"BD"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"2D", X"2D", X"2D"), (X"B3", X"B3", X"B3"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"3C", X"3C", X"3C"), (X"A4", X"A4", X"A4"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"02", X"02", X"02"), (X"29", X"29", X"29"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"32", X"32", X"32"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"93", X"93", X"93"), (X"4A", X"4A", X"4A"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"A2", X"A2", X"A2"), (X"3B", X"3B", X"3B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"B1", X"B1", X"B1"), (X"2C", X"2C", X"2C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"C5", X"C5", X"C5"), (X"18", X"18", X"18"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"D0", X"D0", X"D0"), (X"0E", X"0E", X"0E"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"D6", X"D6", X"D6"), (X"04", X"04", X"04"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"0D", X"0D", X"0D"), (X"D0", X"D0", X"D0"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"17", X"17", X"17"), (X"C6", X"C6", X"C6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"21", X"21", X"21"), (X"BC", X"BC", X"BC"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2B", X"2B", X"2B"), (X"B2", X"B2", X"B2"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"3A", X"3A", X"3A"), (X"A3", X"A3", X"A3"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2A", X"2A", X"2A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"36", X"36", X"36"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"93", X"93", X"93"), (X"4A", X"4A", X"4A"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"A2", X"A2", X"A2"), (X"3B", X"3B", X"3B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"B1", X"B1", X"B1"), (X"2C", X"2C", X"2C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"C5", X"C5", X"C5"), (X"18", X"18", X"18"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"D0", X"D0", X"D0"), (X"0E", X"0E", X"0E"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"D6", X"D6", X"D6"), (X"04", X"04", X"04"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"0D", X"0D", X"0D"), (X"D0", X"D0", X"D0"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"17", X"17", X"17"), (X"C6", X"C6", X"C6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"21", X"21", X"21"), (X"BC", X"BC", X"BC"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2B", X"2B", X"2B"), (X"B2", X"B2", X"B2"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"3A", X"3A", X"3A"), (X"A3", X"A3", X"A3"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2E", X"2E", X"2E"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"3C", X"3C", X"3C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"93", X"93", X"93"), (X"4A", X"4A", X"4A"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"A2", X"A2", X"A2"), (X"3B", X"3B", X"3B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"B1", X"B1", X"B1"), (X"2C", X"2C", X"2C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"C5", X"C5", X"C5"), (X"18", X"18", X"18"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"D0", X"D0", X"D0"), (X"0E", X"0E", X"0E"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"D6", X"D6", X"D6"), (X"04", X"04", X"04"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"0D", X"0D", X"0D"), (X"D0", X"D0", X"D0"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"17", X"17", X"17"), (X"C6", X"C6", X"C6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"21", X"21", X"21"), (X"BC", X"BC", X"BC"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2B", X"2B", X"2B"), (X"B2", X"B2", X"B2"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"3A", X"3A", X"3A"), (X"A3", X"A3", X"A3"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"34", X"34", X"34"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"0B", X"0B", X"0B"), (X"0B", X"0B", X"0B"), (X"0B", X"0B", X"0B"), (X"0B", X"0B", X"0B"), (X"0B", X"0B", X"0B"), (X"0B", X"0B", X"0B"), (X"6D", X"6D", X"6D"), (X"BE", X"BA", X"BB"), (X"85", X"7D", X"7F"), (X"85", X"7D", X"7F"), (X"85", X"7D", X"7F"), (X"85", X"7D", X"7F"), (X"85", X"7D", X"7F"), (X"85", X"7D", X"7F"), (X"85", X"7D", X"7F"), (X"85", X"7D", X"7F"), (X"85", X"7D", X"7F"), (X"BD", X"B9", X"BA"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"AC", X"AC", X"AC"), (X"7F", X"7F", X"7F"), (X"7F", X"7F", X"7F"), (X"7F", X"7F", X"7F"), (X"7F", X"7F", X"7F"), (X"47", X"47", X"47"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"93", X"93", X"93"), (X"4A", X"4A", X"4A"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"A2", X"A2", X"A2"), (X"3B", X"3B", X"3B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"B1", X"B1", X"B1"), (X"2C", X"2C", X"2C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"C5", X"C5", X"C5"), (X"18", X"18", X"18"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"D0", X"D0", X"D0"), (X"0E", X"0E", X"0E"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"D6", X"D6", X"D6"), (X"04", X"04", X"04"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"0D", X"0D", X"0D"), (X"D0", X"D0", X"D0"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"17", X"17", X"17"), (X"C6", X"C6", X"C6"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"21", X"21", X"21"), (X"BC", X"BC", X"BC"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2B", X"2B", X"2B"), (X"B2", X"B2", X"B2"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"3A", X"3A", X"3A"), (X"A3", X"A3", X"A3"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"3F", X"3F", X"3F"), (X"7F", X"7F", X"7F"), (X"7F", X"7F", X"7F"), (X"7F", X"7F", X"7F"), (X"7F", X"7F", X"7F"), (X"A4", X"A4", X"A4"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"C2", X"C1", X"C6"), (X"7F", X"7E", X"89"), (X"7F", X"7E", X"89"), (X"7F", X"7E", X"89"), (X"7F", X"7E", X"89"), (X"7F", X"7E", X"89"), (X"7F", X"7E", X"89"), (X"7F", X"7E", X"89"), (X"7F", X"7E", X"89"), (X"7F", X"7E", X"89"), (X"B3", X"B2", X"B9"), (X"7C", X"7C", X"7C"), (X"0B", X"0B", X"0B"), (X"0B", X"0B", X"0B"), (X"0B", X"0B", X"0B"), (X"0B", X"0B", X"0B"), (X"0B", X"0B", X"0B"), (X"0B", X"0B", X"0B"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"DA", X"DA", X"DA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"DA", X"DA", X"DA"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"D2", X"D2", X"D2"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"75", X"75", X"75"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"20", X"20", X"20"), (X"10", X"10", X"10"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"39", X"39", X"39"), (X"AD", X"AD", X"AD"), (X"AD", X"AD", X"AD"), (X"41", X"41", X"41"), (X"08", X"08", X"08"), (X"7B", X"7B", X"7B"), (X"C5", X"C5", X"C5"), (X"9C", X"9C", X"9C"), (X"2D", X"2D", X"2D"), (X"0E", X"0E", X"0E"), (X"6D", X"6D", X"6D"), (X"BF", X"BF", X"BF"), (X"88", X"88", X"88"), (X"1C", X"1C", X"1C"), (X"19", X"19", X"19"), (X"84", X"84", X"84"), (X"E7", X"E7", X"E7"), (X"7C", X"7C", X"7C"), (X"10", X"10", X"10"), (X"29", X"29", X"29"), (X"98", X"98", X"98"), (X"BB", X"BB", X"BB"), (X"35", X"35", X"35"), (X"88", X"88", X"88"), (X"4C", X"4C", X"4C"), (X"6E", X"6E", X"6E"), (X"66", X"66", X"66"), (X"7D", X"7D", X"7D"), (X"88", X"88", X"88"), (X"3B", X"3B", X"3B"), (X"95", X"95", X"95"), (X"2C", X"2C", X"2C"), (X"A1", X"A1", X"A1"), (X"24", X"24", X"24"), (X"A5", X"A5", X"A5"), (X"23", X"23", X"23"), (X"9F", X"9F", X"9F"), (X"31", X"31", X"31"), (X"B7", X"B7", X"B7"), (X"4C", X"4C", X"4C"), (X"75", X"75", X"75"), (X"5F", X"5F", X"5F"), (X"5B", X"5B", X"5B"), (X"78", X"78", X"78"), (X"6E", X"6E", X"6E"), (X"47", X"47", X"47"), (X"62", X"62", X"62"), (X"84", X"84", X"84"), (X"5B", X"5B", X"5B"), (X"6D", X"6D", X"6D"), (X"09", X"09", X"09"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"67", X"67", X"67"), (X"72", X"72", X"72"), (X"7C", X"7C", X"7C"), (X"50", X"50", X"50"), (X"50", X"50", X"50"), (X"7F", X"7F", X"7F"), (X"63", X"63", X"63"), (X"64", X"64", X"64"), (X"65", X"65", X"65"), (X"65", X"65", X"65"), (X"69", X"69", X"69"), (X"93", X"93", X"93"), (X"65", X"65", X"65"), (X"62", X"62", X"62"), (X"63", X"63", X"63"), (X"64", X"64", X"64"), (X"65", X"65", X"65"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"62", X"62", X"62"), (X"62", X"62", X"62"), (X"68", X"68", X"68"), (X"90", X"90", X"90"), (X"65", X"65", X"65"), (X"66", X"66", X"66"), (X"62", X"62", X"62"), (X"61", X"61", X"61"), (X"5C", X"5C", X"5C"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"70", X"70", X"70"), (X"6E", X"6E", X"6E"), (X"5A", X"5A", X"5A"), (X"89", X"89", X"89"), (X"6C", X"6C", X"6C"), (X"6D", X"6D", X"6D"), (X"59", X"59", X"59"), (X"56", X"56", X"56"), (X"74", X"74", X"74"), (X"69", X"69", X"69"), (X"5B", X"5B", X"5B"), (X"5A", X"5A", X"5A"), (X"6C", X"6C", X"6C"), (X"7D", X"7D", X"7D"), (X"7A", X"7A", X"7A"), (X"5D", X"5D", X"5D"), (X"6D", X"6D", X"6D"), (X"6D", X"6D", X"6D"), (X"5D", X"5D", X"5D"), (X"4F", X"4F", X"4F"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"0D", X"0D", X"0D"), (X"24", X"24", X"24"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"6A", X"6A", X"6A"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"CE", X"CE", X"CE"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"DE", X"DE", X"DE"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"D6", X"D6", X"D6"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"5A", X"5A", X"5A"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"52", X"52", X"52"), (X"08", X"08", X"08"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"02", X"02"), (X"48", X"48", X"48"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"52", X"52", X"52"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"67", X"67", X"67"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"52", X"52", X"52"), (X"08", X"08", X"08"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"02", X"02"), (X"48", X"48", X"48"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"60", X"60", X"60"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"72", X"72", X"72"), (X"05", X"05", X"05"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"52", X"52", X"52"), (X"08", X"08", X"08"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"02", X"02"), (X"48", X"48", X"48"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"6C", X"6C", X"6C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"78", X"78", X"78"), (X"10", X"10", X"10"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"52", X"52", X"52"), (X"08", X"08", X"08"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"02", X"02"), (X"48", X"48", X"48"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"0A", X"0A", X"0A"), (X"76", X"76", X"76"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"52", X"52", X"52"), (X"08", X"08", X"08"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"02", X"02"), (X"48", X"48", X"48"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"1A", X"1A", X"1A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"37", X"37", X"37"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"52", X"52", X"52"), (X"08", X"08", X"08"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"02", X"02"), (X"48", X"48", X"48"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2F", X"2F", X"2F"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B7", X"B9", X"B8"), (X"78", X"7B", X"7A"), (X"78", X"7B", X"7A"), (X"78", X"7B", X"7A"), (X"78", X"7B", X"7A"), (X"78", X"7B", X"7A"), (X"78", X"7B", X"7A"), (X"78", X"7B", X"7A"), (X"78", X"7B", X"7A"), (X"78", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"4E", X"4E", X"4E"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"52", X"52", X"52"), (X"08", X"08", X"08"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"02", X"02"), (X"48", X"48", X"48"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"46", X"46", X"46"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BE"), (X"7A", X"7B", X"77"), (X"7A", X"7B", X"77"), (X"7A", X"7B", X"77"), (X"7A", X"7B", X"77"), (X"7A", X"7B", X"77"), (X"7A", X"7B", X"77"), (X"7A", X"7B", X"77"), (X"7A", X"7B", X"77"), (X"7A", X"7B", X"77"), (X"B0", X"B0", X"AE"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"68", X"68", X"68"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"52", X"52", X"52"), (X"08", X"08", X"08"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"02", X"02"), (X"48", X"48", X"48"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"60", X"60", X"60"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"77", X"77", X"77"), (X"0C", X"0C", X"0C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"52", X"52", X"52"), (X"08", X"08", X"08"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"02", X"02"), (X"48", X"48", X"48"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"08", X"08", X"08"), (X"73", X"73", X"73"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BB", X"C2", X"BF"), (X"7F", X"8C", X"87"), (X"7F", X"8C", X"87"), (X"7F", X"8C", X"87"), (X"7F", X"8C", X"87"), (X"7F", X"8C", X"87"), (X"7F", X"8C", X"87"), (X"7F", X"8C", X"87"), (X"7F", X"8C", X"87"), (X"7F", X"8C", X"87"), (X"BA", X"C1", X"BE"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"B1", X"B1", X"B1"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"2C", X"2C", X"2C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"52", X"52", X"52"), (X"08", X"08", X"08"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"02", X"02", X"02"), (X"48", X"48", X"48"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"23", X"23", X"23"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"A9", X"A9", X"A9"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"C6", X"C7", X"BE"), (X"87", X"8A", X"78"), (X"87", X"8A", X"78"), (X"87", X"8A", X"78"), (X"87", X"8A", X"78"), (X"87", X"8A", X"78"), (X"87", X"8A", X"78"), (X"87", X"8A", X"78"), (X"87", X"8A", X"78"), (X"87", X"8A", X"78"), (X"B8", X"B9", X"AE"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"A6", X"A6", X"A6"), (X"D8", X"D5", X"D6"), (X"B6", X"B0", X"B2"), (X"B6", X"B0", X"B2"), (X"B6", X"B0", X"B2"), (X"B6", X"B0", X"B2"), (X"B6", X"B0", X"B2"), (X"B6", X"B0", X"B2"), (X"B6", X"B0", X"B2"), (X"B6", X"B0", X"B2"), (X"B6", X"B0", X"B2"), (X"D7", X"D4", X"D5"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"CD", X"CD", X"CD"), (X"B2", X"B2", X"B2"), (X"B2", X"B2", X"B2"), (X"B2", X"B2", X"B2"), (X"B2", X"B2", X"B2"), (X"B2", X"B2", X"B2"), (X"B2", X"B2", X"B2"), (X"60", X"60", X"60"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"59", X"59", X"59"), (X"7B", X"7B", X"7B"), (X"84", X"84", X"84"), (X"55", X"55", X"55"), (X"55", X"55", X"55"), (X"9A", X"9A", X"9A"), (X"8A", X"8A", X"8A"), (X"4C", X"4C", X"4C"), (X"68", X"68", X"68"), (X"8C", X"8C", X"8C"), (X"66", X"66", X"66"), (X"55", X"55", X"55"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"55", X"55", X"55"), (X"B2", X"B2", X"B2"), (X"B2", X"B2", X"B2"), (X"B2", X"B2", X"B2"), (X"B2", X"B2", X"B2"), (X"B2", X"B2", X"B2"), (X"B2", X"B2", X"B2"), (X"C8", X"C8", X"C8"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"DA", X"DA", X"DD"), (X"B2", X"B1", X"B8"), (X"B2", X"B1", X"B8"), (X"B2", X"B1", X"B8"), (X"B2", X"B1", X"B8"), (X"B2", X"B1", X"B8"), (X"B2", X"B1", X"B8"), (X"B2", X"B1", X"B8"), (X"B2", X"B1", X"B8"), (X"B2", X"B1", X"B8"), (X"D1", X"D1", X"D5"), (X"B0", X"B0", X"B0"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), (X"6B", X"6B", X"6B"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"66", X"66", X"66"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"5A", X"5A", X"5A"), (X"91", X"91", X"91"), (X"9E", X"9E", X"9E"), (X"64", X"64", X"64"), (X"66", X"66", X"66"), (X"A4", X"A4", X"A4"), (X"8E", X"8E", X"8E"), (X"5B", X"5B", X"5B"), (X"7C", X"7C", X"7C"), (X"A6", X"A6", X"A6"), (X"79", X"79", X"79"), (X"58", X"58", X"58"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"5E", X"5E", X"5E"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"79", X"79", X"79"), (X"10", X"10", X"10"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"5A", X"5A", X"5A"), (X"91", X"91", X"91"), (X"9E", X"9E", X"9E"), (X"64", X"64", X"64"), (X"66", X"66", X"66"), (X"A4", X"A4", X"A4"), (X"8E", X"8E", X"8E"), (X"5B", X"5B", X"5B"), (X"7C", X"7C", X"7C"), (X"A6", X"A6", X"A6"), (X"79", X"79", X"79"), (X"58", X"58", X"58"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"0C", X"0C", X"0C"), (X"76", X"76", X"76"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"36", X"36", X"36"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"5A", X"5A", X"5A"), (X"91", X"91", X"91"), (X"9E", X"9E", X"9E"), (X"64", X"64", X"64"), (X"66", X"66", X"66"), (X"A4", X"A4", X"A4"), (X"8E", X"8E", X"8E"), (X"5B", X"5B", X"5B"), (X"7C", X"7C", X"7C"), (X"A6", X"A6", X"A6"), (X"79", X"79", X"79"), (X"58", X"58", X"58"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2E", X"2E", X"2E"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"5C", X"5C", X"5C"), (X"01", X"01", X"01"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"5A", X"5A", X"5A"), (X"91", X"91", X"91"), (X"9E", X"9E", X"9E"), (X"64", X"64", X"64"), (X"66", X"66", X"66"), (X"A4", X"A4", X"A4"), (X"8E", X"8E", X"8E"), (X"5B", X"5B", X"5B"), (X"7C", X"7C", X"7C"), (X"A6", X"A6", X"A6"), (X"79", X"79", X"79"), (X"58", X"58", X"58"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"55", X"55", X"55"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"78", X"78", X"78"), (X"0F", X"0F", X"0F"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"5A", X"5A", X"5A"), (X"91", X"91", X"91"), (X"9E", X"9E", X"9E"), (X"64", X"64", X"64"), (X"66", X"66", X"66"), (X"A4", X"A4", X"A4"), (X"8E", X"8E", X"8E"), (X"5B", X"5B", X"5B"), (X"7C", X"7C", X"7C"), (X"A6", X"A6", X"A6"), (X"79", X"79", X"79"), (X"58", X"58", X"58"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"0A", X"0A", X"0A"), (X"76", X"76", X"76"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"39", X"39", X"39"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"5A", X"5A", X"5A"), (X"91", X"91", X"91"), (X"9E", X"9E", X"9E"), (X"64", X"64", X"64"), (X"66", X"66", X"66"), (X"A4", X"A4", X"A4"), (X"8E", X"8E", X"8E"), (X"5B", X"5B", X"5B"), (X"7C", X"7C", X"7C"), (X"A6", X"A6", X"A6"), (X"79", X"79", X"79"), (X"58", X"58", X"58"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"31", X"31", X"31"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"65", X"65", X"65"), (X"02", X"02", X"02"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"5A", X"5A", X"5A"), (X"91", X"91", X"91"), (X"9E", X"9E", X"9E"), (X"64", X"64", X"64"), (X"66", X"66", X"66"), (X"A4", X"A4", X"A4"), (X"8E", X"8E", X"8E"), (X"5B", X"5B", X"5B"), (X"7C", X"7C", X"7C"), (X"A6", X"A6", X"A6"), (X"79", X"79", X"79"), (X"58", X"58", X"58"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"5F", X"5F", X"5F"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B8", X"B8", X"B8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B7", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"1F", X"1F", X"1F"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"5A", X"5A", X"5A"), (X"91", X"91", X"91"), (X"9E", X"9E", X"9E"), (X"64", X"64", X"64"), (X"66", X"66", X"66"), (X"A4", X"A4", X"A4"), (X"8E", X"8E", X"8E"), (X"5B", X"5B", X"5B"), (X"7C", X"7C", X"7C"), (X"A6", X"A6", X"A6"), (X"79", X"79", X"79"), (X"58", X"58", X"58"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"18", X"18", X"18"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BF"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"B0", X"B0", X"AF"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"72", X"72", X"72"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"5A", X"5A", X"5A"), (X"91", X"91", X"91"), (X"9E", X"9E", X"9E"), (X"64", X"64", X"64"), (X"66", X"66", X"66"), (X"A4", X"A4", X"A4"), (X"8E", X"8E", X"8E"), (X"5B", X"5B", X"5B"), (X"7C", X"7C", X"7C"), (X"A6", X"A6", X"A6"), (X"79", X"79", X"79"), (X"58", X"58", X"58"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"7F", X"7F", X"7F"), (X"CA", X"C0", X"C3"), (X"9C", X"89", X"8F"), (X"9C", X"89", X"8F"), (X"9C", X"89", X"8F"), (X"9C", X"89", X"8F"), (X"9C", X"89", X"8F"), (X"9C", X"89", X"8F"), (X"9C", X"89", X"8F"), (X"9C", X"89", X"8F"), (X"9C", X"89", X"8F"), (X"CA", X"BF", X"C2"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"B6", X"B6", X"B6"), (X"8F", X"8F", X"8F"), (X"8F", X"8F", X"8F"), (X"8F", X"8F", X"8F"), (X"8F", X"8F", X"8F"), (X"8F", X"8F", X"8F"), (X"8F", X"8F", X"8F"), (X"8F", X"8F", X"8F"), (X"8F", X"8F", X"8F"), (X"8F", X"8F", X"8F"), (X"C6", X"C6", X"C6"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"DD", X"DD", X"DD"), (X"DD", X"DD", X"DD"), (X"53", X"53", X"53"), (X"0A", X"0A", X"0A"), (X"70", X"70", X"70"), (X"EC", X"EC", X"EC"), (X"C8", X"C8", X"C8"), (X"3A", X"3A", X"3A"), (X"12", X"12", X"12"), (X"8C", X"8C", X"8C"), (X"F5", X"F5", X"F5"), (X"AF", X"AF", X"AF"), (X"24", X"24", X"24"), (X"20", X"20", X"20"), (X"A9", X"A9", X"A9"), (X"F6", X"F6", X"F6"), (X"93", X"93", X"93"), (X"14", X"14", X"14"), (X"34", X"34", X"34"), (X"C3", X"C3", X"C3"), (X"EF", X"EF", X"EF"), (X"44", X"44", X"44"), (X"AE", X"AE", X"AE"), (X"61", X"61", X"61"), (X"8D", X"8D", X"8D"), (X"83", X"83", X"83"), (X"6B", X"6B", X"6B"), (X"A5", X"A5", X"A5"), (X"4B", X"4B", X"4B"), (X"BF", X"BF", X"BF"), (X"38", X"38", X"38"), (X"CE", X"CE", X"CE"), (X"2D", X"2D", X"2D"), (X"D4", X"D4", X"D4"), (X"2C", X"2C", X"2C"), (X"CB", X"CB", X"CB"), (X"3F", X"3F", X"3F"), (X"B3", X"B3", X"B3"), (X"5A", X"5A", X"5A"), (X"96", X"96", X"96"), (X"7A", X"7A", X"7A"), (X"75", X"75", X"75"), (X"9A", X"9A", X"9A"), (X"8C", X"8C", X"8C"), (X"5A", X"5A", X"5A"), (X"7D", X"7D", X"7D"), (X"A9", X"A9", X"A9"), (X"75", X"75", X"75"), (X"5A", X"5A", X"5A"), (X"91", X"91", X"91"), (X"9E", X"9E", X"9E"), (X"64", X"64", X"64"), (X"66", X"66", X"66"), (X"A4", X"A4", X"A4"), (X"8E", X"8E", X"8E"), (X"5B", X"5B", X"5B"), (X"7C", X"7C", X"7C"), (X"A6", X"A6", X"A6"), (X"79", X"79", X"79"), (X"58", X"58", X"58"), (X"92", X"92", X"92"), (X"9F", X"9F", X"9F"), (X"66", X"66", X"66"), (X"67", X"67", X"67"), (X"A2", X"A2", X"A2"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"81", X"81", X"81"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"80", X"80", X"80"), (X"82", X"82", X"82"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7D", X"7D", X"7D"), (X"7E", X"7E", X"7E"), (X"7F", X"7F", X"7F"), (X"81", X"81", X"81"), (X"82", X"82", X"82"), (X"83", X"83", X"83"), (X"7E", X"7E", X"7E"), (X"7D", X"7D", X"7D"), (X"76", X"76", X"76"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"90", X"90", X"90"), (X"8D", X"8D", X"8D"), (X"6A", X"6A", X"6A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"72", X"72", X"72"), (X"6E", X"6E", X"6E"), (X"95", X"95", X"95"), (X"86", X"86", X"86"), (X"74", X"74", X"74"), (X"74", X"74", X"74"), (X"8A", X"8A", X"8A"), (X"94", X"94", X"94"), (X"6A", X"6A", X"6A"), (X"77", X"77", X"77"), (X"8B", X"8B", X"8B"), (X"8B", X"8B", X"8B"), (X"77", X"77", X"77"), (X"65", X"65", X"65"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"16", X"16", X"16"), (X"C9", X"C9", X"C9"), (X"8F", X"8F", X"8F"), (X"8F", X"8F", X"8F"), (X"8F", X"8F", X"8F"), (X"8F", X"8F", X"8F"), (X"8F", X"8F", X"8F"), (X"8F", X"8F", X"8F"), (X"8F", X"8F", X"8F"), (X"8F", X"8F", X"8F"), (X"8F", X"8F", X"8F"), (X"AF", X"AF", X"AF"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"C9", X"C7", X"D4"), (X"8F", X"8B", X"A6"), (X"8F", X"8B", X"A6"), (X"8F", X"8B", X"A6"), (X"8F", X"8B", X"A6"), (X"8F", X"8B", X"A6"), (X"8F", X"8B", X"A6"), (X"8F", X"8B", X"A6"), (X"8F", X"8B", X"A6"), (X"8F", X"8B", X"A6"), (X"BC", X"BA", X"CA"), (X"8C", X"8C", X"8C"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"CE", X"D4", X"D2"), (X"A3", X"AE", X"AA"), (X"A3", X"AE", X"AA"), (X"A3", X"AE", X"AA"), (X"A3", X"AE", X"AA"), (X"A3", X"AE", X"AA"), (X"A3", X"AE", X"AA"), (X"A3", X"AE", X"AA"), (X"A3", X"AE", X"AA"), (X"A3", X"AE", X"AA"), (X"CD", X"D3", X"D1"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"C8", X"C8", X"C8"), (X"AA", X"AA", X"AA"), (X"AA", X"AA", X"AA"), (X"AA", X"AA", X"AA"), (X"AA", X"AA", X"AA"), (X"AA", X"AA", X"AA"), (X"AA", X"AA", X"AA"), (X"AA", X"AA", X"AA"), (X"AA", X"AA", X"AA"), (X"AA", X"AA", X"AA"), (X"DB", X"DB", X"DB"), (X"70", X"70", X"70"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"07", X"07", X"07"), (X"16", X"16", X"16"), (X"16", X"16", X"16"), (X"08", X"08", X"08"), (X"01", X"01", X"01"), (X"0B", X"0B", X"0B"), (X"18", X"18", X"18"), (X"14", X"14", X"14"), (X"06", X"06", X"06"), (X"02", X"02", X"02"), (X"0E", X"0E", X"0E"), (X"3A", X"3A", X"3A"), (X"40", X"40", X"40"), (X"32", X"32", X"32"), (X"31", X"31", X"31"), (X"3F", X"3F", X"3F"), (X"47", X"47", X"47"), (X"3D", X"3D", X"3D"), (X"30", X"30", X"30"), (X"33", X"33", X"33"), (X"41", X"41", X"41"), (X"46", X"46", X"46"), (X"35", X"35", X"35"), (X"3F", X"3F", X"3F"), (X"38", X"38", X"38"), (X"3C", X"3C", X"3C"), (X"3B", X"3B", X"3B"), (X"39", X"39", X"39"), (X"3F", X"3F", X"3F"), (X"35", X"35", X"35"), (X"41", X"41", X"41"), (X"34", X"34", X"34"), (X"43", X"43", X"43"), (X"5A", X"5A", X"5A"), (X"71", X"71", X"71"), (X"60", X"60", X"60"), (X"70", X"70", X"70"), (X"62", X"62", X"62"), (X"6E", X"6E", X"6E"), (X"65", X"65", X"65"), (X"6B", X"6B", X"6B"), (X"68", X"68", X"68"), (X"68", X"68", X"68"), (X"6B", X"6B", X"6B"), (X"6A", X"6A", X"6A"), (X"65", X"65", X"65"), (X"68", X"68", X"68"), (X"6D", X"6D", X"6D"), (X"67", X"67", X"67"), (X"64", X"64", X"64"), (X"6A", X"6A", X"6A"), (X"6B", X"6B", X"6B"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"6C", X"6C", X"6C"), (X"97", X"97", X"97"), (X"93", X"93", X"93"), (X"96", X"96", X"96"), (X"9A", X"9A", X"9A"), (X"96", X"96", X"96"), (X"92", X"92", X"92"), (X"98", X"98", X"98"), (X"99", X"99", X"99"), (X"94", X"94", X"94"), (X"94", X"94", X"94"), (X"9A", X"9A", X"9A"), (X"96", X"96", X"96"), (X"96", X"96", X"96"), (X"97", X"97", X"97"), (X"97", X"97", X"97"), (X"97", X"97", X"97"), (X"97", X"97", X"97"), (X"97", X"97", X"97"), (X"96", X"96", X"96"), (X"96", X"96", X"96"), (X"96", X"96", X"96"), (X"9B", X"9B", X"9B"), (X"C4", X"C4", X"C4"), (X"C4", X"C4", X"C4"), (X"C4", X"C4", X"C4"), (X"C4", X"C4", X"C4"), (X"C4", X"C4", X"C4"), (X"C4", X"C4", X"C4"), (X"C5", X"C5", X"C5"), (X"C5", X"C5", X"C5"), (X"C4", X"C4", X"C4"), (X"C4", X"C4", X"C4"), (X"C3", X"C3", X"C3"), (X"C3", X"C3", X"C3"), (X"C3", X"C3", X"C3"), (X"C6", X"C6", X"C6"), (X"C6", X"C6", X"C6"), (X"C2", X"C2", X"C2"), (X"C4", X"C4", X"C4"), (X"C5", X"C5", X"C5"), (X"C5", X"C5", X"C5"), (X"C3", X"C3", X"C3"), (X"C2", X"C2", X"C2"), (X"D0", X"D0", X"D0"), (X"F3", X"F3", X"F3"), (X"F1", X"F1", X"F1"), (X"F1", X"F1", X"F1"), (X"F3", X"F3", X"F3"), (X"F4", X"F4", X"F4"), (X"F0", X"F0", X"F0"), (X"F1", X"F1", X"F1"), (X"F3", X"F3", X"F3"), (X"F3", X"F3", X"F3"), (X"F1", X"F1", X"F1"), (X"F0", X"F0", X"F0"), (X"E5", X"E5", X"E5"), (X"E5", X"E5", X"E5"), (X"E5", X"E5", X"E5"), (X"E5", X"E5", X"E5"), (X"CD", X"CD", X"CD"), (X"E0", X"E0", X"E0"), (X"AA", X"AA", X"AA"), (X"AA", X"AA", X"AA"), (X"AA", X"AA", X"AA"), (X"AA", X"AA", X"AA"), (X"AA", X"AA", X"AA"), (X"AA", X"AA", X"AA"), (X"AA", X"AA", X"AA"), (X"AA", X"AA", X"AA"), (X"AA", X"AA", X"AA"), (X"C2", X"C2", X"C2"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"D6", X"D8", X"D0"), (X"AA", X"AD", X"9D"), (X"AA", X"AD", X"9D"), (X"AA", X"AD", X"9D"), (X"AA", X"AD", X"9D"), (X"AA", X"AD", X"9D"), (X"AA", X"AD", X"9D"), (X"AA", X"AD", X"9D"), (X"AA", X"AD", X"9D"), (X"AA", X"AD", X"9D"), (X"CC", X"CE", X"C5"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"99", X"99", X"99"), (X"0C", X"0C", X"0C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"5E", X"5E", X"5E"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"97", X"97", X"97"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"9D", X"9D", X"9D"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"D6", X"D6", X"D6"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F6", X"F6", X"F6"), (X"A4", X"A4", X"A4"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"41", X"41", X"41"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"5E", X"5E", X"5E"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"97", X"97", X"97"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"9D", X"9D", X"9D"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"D6", X"D6", X"D6"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"C0", X"C0", X"C0"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"73", X"73", X"73"), (X"0D", X"0D", X"0D"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"5E", X"5E", X"5E"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"97", X"97", X"97"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"9D", X"9D", X"9D"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"D6", X"D6", X"D6"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F5", X"F5", X"F5"), (X"86", X"86", X"86"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"49", X"49", X"49"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"5E", X"5E", X"5E"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"97", X"97", X"97"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"9D", X"9D", X"9D"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"D6", X"D6", X"D6"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B7", X"B7", X"B7"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"78", X"78", X"78"), (X"16", X"16", X"16"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"5E", X"5E", X"5E"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"97", X"97", X"97"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"9D", X"9D", X"9D"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"D6", X"D6", X"D6"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"EC", X"EC", X"EC"), (X"80", X"80", X"80"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"5A", X"5A", X"5A"), (X"01", X"01", X"01"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"5E", X"5E", X"5E"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"97", X"97", X"97"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"9D", X"9D", X"9D"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"D6", X"D6", X"D6"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"A4", X"A4", X"A4"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"2C", X"2C", X"2C"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"5E", X"5E", X"5E"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"97", X"97", X"97"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"9D", X"9D", X"9D"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"D6", X"D6", X"D6"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"D6", X"D6", X"D6"), (X"7B", X"7B", X"7B"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"6F", X"6F", X"6F"), (X"0B", X"0B", X"0B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"5E", X"5E", X"5E"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"97", X"97", X"97"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"9D", X"9D", X"9D"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"D6", X"D6", X"D6"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F8", X"F8", X"F8"), (X"8A", X"8A", X"8A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"50", X"50", X"50"), (X"01", X"01", X"01"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"5E", X"5E", X"5E"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"97", X"97", X"97"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"9D", X"9D", X"9D"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"D6", X"D6", X"D6"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"DD", X"B0", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"76", X"76", X"76"), (X"1B", X"1B", X"1B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"33", X"33", X"33"), (X"5E", X"5E", X"5E"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"66", X"66", X"66"), (X"97", X"97", X"97"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"99", X"99", X"99"), (X"9D", X"9D", X"9D"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"CC", X"CC", X"CC"), (X"D6", X"D6", X"D6"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"E8", X"E8", X"E8"), (X"7F", X"7F", X"7F"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"BE", X"F6"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"B7", X"B7", X"B7"), (X"DC", X"DE", X"DD"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"BD", X"C1", X"BF"), (X"DB", X"DD", X"DC"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"CB", X"88", X"9B"), (X"D0", X"C0", X"94"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"EB", X"E4", X"D2"), (X"D1", X"D1", X"D1"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"A9", X"A9", X"A9"), (X"B2", X"B2", X"B2"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"BA", X"BA", X"BA"), (X"C4", X"C4", X"C4"), (X"C8", X"C8", X"C8"), (X"C8", X"C8", X"C8"), (X"C8", X"C8", X"C8"), (X"C8", X"C8", X"C8"), (X"C8", X"C8", X"C8"), (X"C8", X"C8", X"C8"), (X"C8", X"C8", X"C8"), (X"C8", X"C8", X"C8"), (X"C8", X"C8", X"C8"), (X"C8", X"C8", X"C8"), (X"35", X"35", X"35"), (X"0E", X"0E", X"0E"), (X"0E", X"0E", X"0E"), (X"0E", X"0E", X"0E"), (X"0E", X"0E", X"0E"), (X"97", X"97", X"97"), (X"27", X"27", X"27"), (X"0E", X"0E", X"0E"), (X"0E", X"0E", X"0E"), (X"0E", X"0E", X"0E"), (X"0E", X"0E", X"0E"), (X"1A", X"1A", X"1A"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"1C", X"1C", X"1C"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"29", X"29", X"29"), (X"2A", X"2A", X"2A"), (X"37", X"37", X"37"), (X"37", X"37", X"37"), (X"37", X"37", X"37"), (X"37", X"37", X"37"), (X"37", X"37", X"37"), (X"37", X"37", X"37"), (X"37", X"37", X"37"), (X"37", X"37", X"37"), (X"37", X"37", X"37"), (X"37", X"37", X"37"), (X"52", X"52", X"52"), (X"F1", X"F1", X"F1"), (X"F1", X"F1", X"F1"), (X"F1", X"F1", X"F1"), (X"F1", X"F1", X"F1"), (X"F1", X"F1", X"F1"), (X"F1", X"F1", X"F1"), (X"F1", X"F1", X"F1"), (X"F1", X"F1", X"F1"), (X"F1", X"F1", X"F1"), (X"F1", X"F1", X"F1"), (X"F4", X"F4", X"F4"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F9", X"F9", X"F9"), (X"C3", X"C3", X"C3"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"BF", X"BF", X"BF"), (X"CD", X"CD", X"CD"), (X"EE", X"E8", X"D8"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"D0", X"BF", X"94"), (X"A6", X"95", X"E2"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"E0", X"E1", X"DE"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"BF", X"C0", X"BB"), (X"D9", X"DA", X"D6"), (X"BF", X"BF", X"BF"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), (X"87", X"87", X"87"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"AA", X"AA", X"AA"), (X"FE", X"FE", X"FE"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"35", X"35", X"35"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FE", X"FE", X"FE"), (X"B2", X"B2", X"B2"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7B", X"7B", X"7B"), (X"C7", X"C7", X"C7"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"35", X"35", X"35"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"CF", X"CF", X"CF"), (X"7B", X"7B", X"7B"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7E", X"7E", X"7E"), (X"DE", X"DE", X"DE"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"35", X"35", X"35"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"E4", X"E4", X"E4"), (X"81", X"81", X"81"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"EF", X"EF", X"EF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"35", X"35", X"35"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F3", X"F3", X"F3"), (X"8B", X"8B", X"8B"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"FD", X"FD", X"FD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"35", X"35", X"35"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FD", X"FD", X"FD"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"76"), (X"7A", X"7B", X"76"), (X"7A", X"7B", X"76"), (X"7A", X"7B", X"76"), (X"7A", X"7B", X"76"), (X"7A", X"7B", X"76"), (X"7A", X"7B", X"76"), (X"7A", X"7B", X"76"), (X"7A", X"7B", X"76"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"B7", X"B7", X"B7"), (X"F7", X"F7", X"F7"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"35", X"35", X"35"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FA", X"FA", X"FA"), (X"B4", X"B4", X"B4"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"9F", X"9F", X"9F"), (X"F9", X"F9", X"F9"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"35", X"35", X"35"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FB", X"FB", X"FB"), (X"A5", X"A5", X"A5"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"A1", X"A1", X"A1"), (X"F9", X"F9", X"F9"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"35", X"35", X"35"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FA", X"FA", X"FA"), (X"A7", X"A7", X"A7"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"9F", X"9F", X"9F"), (X"F7", X"F7", X"F7"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"35", X"35", X"35"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F9", X"F9", X"F9"), (X"A5", X"A5", X"A5"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"0D", X"0D", X"0D"), (X"0D", X"0D", X"0D"), (X"0D", X"0D", X"0D"), (X"0D", X"0D", X"0D"), (X"0D", X"0D", X"0D"), (X"0D", X"0D", X"0D"), (X"6E", X"6E", X"6E"), (X"BF", X"BA", X"BC"), (X"86", X"7E", X"81"), (X"86", X"7E", X"81"), (X"86", X"7E", X"81"), (X"86", X"7E", X"81"), (X"86", X"7E", X"81"), (X"86", X"7E", X"81"), (X"86", X"7E", X"81"), (X"86", X"7E", X"81"), (X"86", X"7E", X"81"), (X"BE", X"B9", X"BB"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A5", X"A5", X"A5"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"D1", X"D1", X"D1"), (X"9E", X"9E", X"9E"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"9F", X"9F", X"9F"), (X"F8", X"F8", X"F8"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"35", X"35", X"35"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"BB", X"BB", X"BB"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"25", X"25", X"25"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F9", X"F9", X"F9"), (X"A5", X"A5", X"A5"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"96", X"96", X"96"), (X"D9", X"D9", X"D9"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"81", X"81", X"81"), (X"9D", X"9D", X"9D"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"C3", X"C2", X"C7"), (X"81", X"7F", X"8B"), (X"81", X"7F", X"8B"), (X"81", X"7F", X"8B"), (X"81", X"7F", X"8B"), (X"81", X"7F", X"8B"), (X"81", X"7F", X"8B"), (X"81", X"7F", X"8B"), (X"81", X"7F", X"8B"), (X"81", X"7F", X"8B"), (X"B4", X"B3", X"BA"), (X"7D", X"7D", X"7D"), (X"0D", X"0D", X"0D"), (X"0D", X"0D", X"0D"), (X"0D", X"0D", X"0D"), (X"0D", X"0D", X"0D"), (X"0D", X"0D", X"0D"), (X"0D", X"0D", X"0D"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"D9", X"DA", X"DA"), (X"B8", X"B9", X"B9"), (X"B8", X"B9", X"B9"), (X"B8", X"B9", X"B9"), (X"B8", X"B9", X"B9"), (X"B8", X"B9", X"B9"), (X"B8", X"B9", X"B9"), (X"B8", X"B9", X"B9"), (X"B8", X"B9", X"B9"), (X"B8", X"B9", X"B9"), (X"D9", X"D9", X"D9"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"CD", X"CD", X"CD"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"E5", X"E5", X"E5"), (X"C9", X"C9", X"C9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B5", X"B5", X"AB"), (X"C3", X"C3", X"46"), (X"CC", X"CC", X"36"), (X"CC", X"CC", X"36"), (X"CC", X"CC", X"36"), (X"CC", X"CC", X"36"), (X"CC", X"CC", X"36"), (X"CC", X"CC", X"36"), (X"CC", X"CC", X"36"), (X"CC", X"CC", X"36"), (X"CC", X"CC", X"36"), (X"A2", X"A2", X"0B"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"BE", X"BE", X"28"), (X"9E", X"9E", X"07"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"8E", X"00"), (X"97", X"08", X"00"), (X"97", X"00", X"00"), (X"97", X"00", X"00"), (X"97", X"00", X"00"), (X"97", X"00", X"00"), (X"97", X"00", X"00"), (X"97", X"00", X"00"), (X"97", X"00", X"00"), (X"97", X"00", X"00"), (X"97", X"02", X"00"), (X"97", X"8B", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"97", X"97", X"00"), (X"9F", X"9F", X"08"), (X"CC", X"CC", X"36"), (X"CC", X"CC", X"36"), (X"CC", X"CC", X"36"), (X"CC", X"CC", X"36"), (X"CC", X"CC", X"36"), (X"CC", X"CC", X"36"), (X"CC", X"CC", X"36"), (X"CC", X"CC", X"36"), (X"CC", X"CC", X"36"), (X"C5", X"C5", X"42"), (X"B5", X"B5", X"A7"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"C5", X"C5", X"C5"), (X"EA", X"EA", X"EA"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"B9", X"B9", X"B9"), (X"C9", X"C9", X"C9"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"DD", X"DE", X"DD"), (X"B9", X"B9", X"B8"), (X"B9", X"B9", X"B8"), (X"B9", X"B9", X"B8"), (X"B9", X"B9", X"B8"), (X"B9", X"B9", X"B8"), (X"B9", X"B9", X"B8"), (X"B9", X"B9", X"B8"), (X"B9", X"B9", X"B8"), (X"B9", X"B9", X"B8"), (X"D5", X"D5", X"D5"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"80", X"80", X"6F"), (X"AE", X"AE", X"1E"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"B4", X"00"), (X"BF", X"0A", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"02", X"00"), (X"BF", X"B0", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"B1", X"B1", X"19"), (X"82", X"82", X"6D"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7C", X"7C", X"76"), (X"A2", X"A2", X"34"), (X"BF", X"BF", X"01"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"B4", X"00"), (X"BF", X"0A", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"02", X"00"), (X"BF", X"B0", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"A5", X"A5", X"2E"), (X"7D", X"7D", X"74"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"79"), (X"92", X"92", X"4E"), (X"BC", X"BC", X"09"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"B4", X"00"), (X"BF", X"0A", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"02", X"00"), (X"BF", X"B0", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BD", X"BD", X"07"), (X"96", X"96", X"48"), (X"7B", X"7B", X"79"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CD", X"CD", X"B0"), (X"BA", X"BA", X"24"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"B4", X"00"), (X"BF", X"0A", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"02", X"00"), (X"BF", X"B0", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"B9", X"B9", X"1E"), (X"D2", X"D2", X"AE"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"93", X"93", X"8D"), (X"9C", X"9C", X"3E"), (X"BC", X"BC", X"04"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"B4", X"00"), (X"BF", X"0A", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"02", X"00"), (X"BF", X"B0", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BD", X"BD", X"03"), (X"9F", X"9F", X"39"), (X"8E", X"8E", X"86"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BA", X"B8", X"B8"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"7D", X"79", X"7A"), (X"B9", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"64"), (X"AF", X"AF", X"1C"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"B4", X"00"), (X"BF", X"0A", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"02", X"00"), (X"BF", X"B0", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"B2", X"B2", X"18"), (X"88", X"88", X"60"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"BF", X"C2"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"7A", X"79", X"7F"), (X"B0", X"AF", X"B3"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B8", X"B8", X"B8"), (X"79", X"7A", X"7A"), (X"79", X"7A", X"7A"), (X"79", X"7A", X"7A"), (X"79", X"7A", X"7A"), (X"79", X"7A", X"7A"), (X"79", X"7A", X"7A"), (X"79", X"7A", X"7A"), (X"79", X"7A", X"7A"), (X"79", X"7A", X"7A"), (X"B7", X"B7", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7B", X"7B", X"79"), (X"94", X"94", X"4B"), (X"B9", X"B9", X"0A"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"B4", X"00"), (X"BF", X"0A", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"02", X"00"), (X"BF", X"B0", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BA", X"BA", X"09"), (X"97", X"97", X"46"), (X"7B", X"7B", X"78"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BF"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"7A", X"7A", X"79"), (X"B0", X"B0", X"AF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7E", X"7E", X"72"), (X"9F", X"9F", X"39"), (X"BC", X"BC", X"06"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"B4", X"00"), (X"BF", X"0A", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"02", X"00"), (X"BF", X"B0", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BC", X"BC", X"04"), (X"A1", X"A1", X"35"), (X"80", X"80", X"70"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"D5", X"9D", X"B0"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B8", X"5A", X"7A"), (X"B6", X"5D", X"72"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"D6", X"C7", X"A0"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"82", X"82", X"6C"), (X"A3", X"A3", X"32"), (X"BC", X"BC", X"05"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"B4", X"00"), (X"BF", X"0A", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"02", X"00"), (X"BF", X"B0", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BD", X"BD", X"04"), (X"A5", X"A5", X"2E"), (X"84", X"84", X"69"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"DC", X"CF", X"AE"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"9D", X"7A", X"1E"), (X"7F", X"67", X"CB"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"7A", X"64", X"E9"), (X"A8", X"9A", X"F0"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"BB", X"C2", X"C0"), (X"7F", X"8D", X"88"), (X"7F", X"8D", X"88"), (X"7F", X"8D", X"88"), (X"7F", X"8D", X"88"), (X"7F", X"8D", X"88"), (X"7F", X"8D", X"88"), (X"7F", X"8D", X"88"), (X"7F", X"8D", X"88"), (X"7F", X"8D", X"88"), (X"BA", X"C1", X"BF"), (X"DA", X"A8", X"B9"), (X"C0", X"6C", X"88"), (X"C0", X"6C", X"88"), (X"C0", X"6C", X"88"), (X"C0", X"6C", X"88"), (X"C0", X"6C", X"88"), (X"C0", X"6C", X"88"), (X"C0", X"6C", X"88"), (X"C0", X"6C", X"88"), (X"C0", X"6C", X"88"), (X"BE", X"6E", X"81"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"DA", X"CD", X"AA"), (X"AA", X"AA", X"AA"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"D4", X"D4", X"D4"), (X"A3", X"A3", X"A3"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"DB", X"DB", X"DB"), (X"9C", X"9C", X"9C"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"91", X"91", X"79"), (X"CC", X"CC", X"63"), (X"C3", X"C3", X"0F"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"B4", X"00"), (X"BF", X"0A", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"02", X"00"), (X"BF", X"B0", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"C2", X"C2", X"0E"), (X"CE", X"CE", X"5F"), (X"92", X"92", X"77"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"98", X"98", X"98"), (X"E0", X"E0", X"E0"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"9C", X"9C", X"9C"), (X"DB", X"DB", X"DB"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"88", X"88", X"88"), (X"A3", X"A3", X"A3"), (X"E0", X"D4", X"B7"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"A8", X"88", X"36"), (X"8D", X"78", X"D0"), (X"88", X"75", X"EB"), (X"88", X"75", X"EB"), (X"88", X"75", X"EB"), (X"88", X"75", X"EB"), (X"88", X"75", X"EB"), (X"88", X"75", X"EB"), (X"88", X"75", X"EB"), (X"88", X"75", X"EB"), (X"88", X"75", X"EB"), (X"B1", X"A5", X"F2"), (X"C6", X"C8", X"BE"), (X"88", X"8C", X"78"), (X"88", X"8C", X"78"), (X"88", X"8C", X"78"), (X"88", X"8C", X"78"), (X"88", X"8C", X"78"), (X"88", X"8C", X"78"), (X"88", X"8C", X"78"), (X"88", X"8C", X"78"), (X"88", X"8C", X"78"), (X"B8", X"BA", X"AE"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"69", X"69", X"69"), (X"69", X"69", X"69"), (X"69", X"69", X"69"), (X"69", X"69", X"69"), (X"69", X"69", X"69"), (X"69", X"69", X"69"), (X"A5", X"A5", X"A5"), (X"D8", X"D4", X"D5"), (X"B5", X"AF", X"B1"), (X"B5", X"AF", X"B1"), (X"B5", X"AF", X"B1"), (X"B5", X"AF", X"B1"), (X"B5", X"AF", X"B1"), (X"B5", X"AF", X"B1"), (X"B5", X"AF", X"B1"), (X"B5", X"AF", X"B1"), (X"B5", X"AF", X"B1"), (X"D7", X"D4", X"D5"), (X"D1", X"D1", X"D1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"D9", X"D9", X"D9"), (X"CC", X"CC", X"CC"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"DE", X"DE", X"DE"), (X"C8", X"C8", X"C8"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"E3", X"E3", X"E3"), (X"C3", X"C3", X"C3"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"E7", X"E7", X"E7"), (X"BE", X"BE", X"BE"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"EA", X"EA", X"EA"), (X"B7", X"B7", X"A9"), (X"9D", X"9D", X"49"), (X"B4", X"B4", X"14"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"B4", X"00"), (X"BF", X"0A", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"02", X"00"), (X"BF", X"B0", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"B5", X"B5", X"12"), (X"9D", X"9D", X"44"), (X"B2", X"B2", X"A1"), (X"EE", X"EE", X"EE"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"BB", X"BB", X"BB"), (X"EB", X"EB", X"EB"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"BE", X"BE", X"BE"), (X"E7", X"E7", X"E7"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"C3", X"C3", X"C3"), (X"E3", X"E3", X"E3"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"C7", X"C7", X"C7"), (X"DE", X"DE", X"DE"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"B1", X"B1", X"B1"), (X"CC", X"CC", X"CC"), (X"DA", X"D9", X"DD"), (X"B1", X"AF", X"B8"), (X"B1", X"AF", X"B8"), (X"B1", X"AF", X"B8"), (X"B1", X"AF", X"B8"), (X"B1", X"AF", X"B8"), (X"B1", X"AF", X"B8"), (X"B1", X"AF", X"B8"), (X"B1", X"AF", X"B8"), (X"B1", X"AF", X"B8"), (X"D1", X"CF", X"D5"), (X"AE", X"AE", X"AE"), (X"69", X"69", X"69"), (X"69", X"69", X"69"), (X"69", X"69", X"69"), (X"69", X"69", X"69"), (X"69", X"69", X"69"), (X"69", X"69", X"69"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"79"), (X"8C", X"8C", X"5A"), (X"A4", X"A4", X"2F"), (X"BB", X"BB", X"07"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"B4", X"00"), (X"BF", X"0A", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"02", X"00"), (X"BF", X"B0", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BC", X"BC", X"05"), (X"A5", X"A5", X"2D"), (X"8D", X"8D", X"57"), (X"7B", X"7B", X"79"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7C", X"7C", X"76"), (X"90", X"90", X"52"), (X"A6", X"A6", X"2C"), (X"BA", X"BA", X"09"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"B4", X"00"), (X"BF", X"0A", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"02", X"00"), (X"BF", X"B0", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BB", X"BB", X"07"), (X"A7", X"A7", X"2A"), (X"92", X"92", X"50"), (X"7D", X"7D", X"74"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7B", X"7B", X"79"), (X"89", X"89", X"5F"), (X"CD", X"CD", X"6E"), (X"B4", X"B4", X"24"), (X"BC", X"BC", X"06"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"B4", X"00"), (X"BF", X"0A", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"02", X"00"), (X"BF", X"B0", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BD", X"BD", X"04"), (X"B3", X"B3", X"1F"), (X"D1", X"D1", X"6E"), (X"8A", X"8A", X"5D"), (X"7B", X"7B", X"78"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B7", X"B9", X"B8"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"77", X"7B", X"7A"), (X"B6", X"B8", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E1", X"E1", X"E1"), (X"86", X"86", X"86"), (X"7D", X"7D", X"75"), (X"89", X"89", X"60"), (X"95", X"95", X"49"), (X"A2", X"A2", X"33"), (X"B1", X"B1", X"18"), (X"B6", X"B6", X"10"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"B4", X"00"), (X"BF", X"0A", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"00", X"00"), (X"BF", X"02", X"00"), (X"BF", X"B0", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"BF", X"BF", X"00"), (X"B7", X"B7", X"0F"), (X"B2", X"B2", X"16"), (X"A2", X"A2", X"33"), (X"97", X"97", X"47"), (X"8A", X"8A", X"5E"), (X"7D", X"7D", X"74"), (X"81", X"81", X"81"), (X"E6", X"E6", X"E6"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"C0", X"BD"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"7A", X"7B", X"75"), (X"B0", X"B0", X"AD"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"BB", X"B6", X"B8"), (X"80", X"77", X"7A"), (X"80", X"77", X"7A"), (X"80", X"77", X"7A"), (X"80", X"77", X"7A"), (X"80", X"77", X"7A"), (X"80", X"77", X"7A"), (X"80", X"77", X"7A"), (X"80", X"77", X"7A"), (X"80", X"77", X"7A"), (X"BA", X"B5", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E1", X"E1", X"E1"), (X"86", X"86", X"86"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7B", X"7B", X"78"), (X"81", X"81", X"6E"), (X"83", X"83", X"6B"), (X"93", X"93", X"4E"), (X"D8", X"D4", X"93"), (X"9A", X"53", X"4F"), (X"A5", X"2F", X"2F"), (X"A5", X"2E", X"2E"), (X"A5", X"2E", X"2E"), (X"A5", X"2E", X"2E"), (X"A5", X"2E", X"2E"), (X"A5", X"2E", X"2E"), (X"A5", X"2E", X"2E"), (X"A5", X"2E", X"2E"), (X"97", X"4B", X"4A"), (X"DA", X"D5", X"95"), (X"94", X"94", X"4F"), (X"84", X"84", X"69"), (X"81", X"81", X"6E"), (X"7C", X"7C", X"77"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"81", X"81", X"81"), (X"E6", X"E6", X"E6"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"BF", X"C5"), (X"7A", X"78", X"85"), (X"7A", X"78", X"85"), (X"7A", X"78", X"85"), (X"7A", X"78", X"85"), (X"7A", X"78", X"85"), (X"7A", X"78", X"85"), (X"7A", X"78", X"85"), (X"7A", X"78", X"85"), (X"7A", X"78", X"85"), (X"B0", X"AF", X"B6"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B8", X"B8", X"B8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B7", X"B7", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E1", X"E1", X"E1"), (X"86", X"86", X"86"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E6", X"E6", X"E6"), (X"81", X"81", X"81"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7C", X"7C", X"7C"), (X"E9", X"E9", X"E9"), (X"7C", X"7C", X"7C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"81", X"81", X"81"), (X"E6", X"E6", X"E6"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"BF", X"BF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B0", X"B0", X"B0"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B8", X"B8", X"B8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B7", X"B7", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E1", X"E1", X"E1"), (X"86", X"86", X"86"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E6", X"E6", X"E6"), (X"81", X"81", X"81"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7C", X"7C", X"7C"), (X"E9", X"E9", X"E9"), (X"7C", X"7C", X"7C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"81", X"81", X"81"), (X"E6", X"E6", X"E6"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"BF", X"BF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B0", X"B0", X"B0"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B8", X"B8", X"B8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B7", X"B7", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E1", X"E1", X"E1"), (X"86", X"86", X"86"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E6", X"E6", X"E6"), (X"81", X"81", X"81"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7C", X"7C", X"7C"), (X"E9", X"E9", X"E9"), (X"7C", X"7C", X"7C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"81", X"81", X"81"), (X"E6", X"E6", X"E6"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"BF", X"BF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B0", X"B0", X"B0"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"66", X"66", X"66"), (X"B8", X"B8", X"B8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B7", X"B7", X"B7"), (X"B0", X"B0", X"B0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"BF", X"BF", X"BF"), (X"A8", X"A8", X"A8"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"C7", X"C7", X"C7"), (X"A0", X"A0", X"A0"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"CF", X"CF", X"CF"), (X"99", X"99", X"99"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"D6", X"D6", X"D6"), (X"91", X"91", X"91"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"DC", X"DC", X"DC"), (X"8C", X"8C", X"8C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E1", X"E1", X"E1"), (X"86", X"86", X"86"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"E6", X"E6", X"E6"), (X"81", X"81", X"81"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7C", X"7C", X"7C"), (X"E9", X"E9", X"E9"), (X"7C", X"7C", X"7C"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"81", X"81", X"81"), (X"E6", X"E6", X"E6"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"86", X"86", X"86"), (X"E1", X"E1", X"E1"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"8B", X"8B", X"8B"), (X"DC", X"DC", X"DC"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"98", X"98", X"98"), (X"CF", X"CF", X"CF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A0", X"A0", X"A0"), (X"C7", X"C7", X"C7"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"A8", X"A8", X"A8"), (X"BF", X"BF", X"BF"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"7A", X"7A", X"7A"), (X"B0", X"B0", X"B0"), (X"76", X"76", X"76"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), 
	(X"2B", X"2B", X"2B"), (X"2B", X"2B", X"2B"), (X"2B", X"2B", X"2B"), (X"2B", X"2B", X"2B"), (X"2B", X"2B", X"2B"), (X"2B", X"2B", X"2B"), (X"80", X"80", X"80"), (X"C4", X"C4", X"C4"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"C3", X"C3", X"C3"), (X"BD", X"BD", X"BD"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"CA", X"CA", X"CA"), (X"B7", X"B7", X"B7"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"D0", X"D0", X"D0"), (X"B0", X"B0", X"B0"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"D7", X"D7", X"D7"), (X"AA", X"AA", X"AA"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"DD", X"DD", X"DD"), (X"A3", X"A3", X"A3"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"E2", X"E2", X"E2"), (X"9F", X"9F", X"9F"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"E6", X"E6", X"E6"), (X"9A", X"9A", X"9A"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"EA", X"EA", X"EA"), (X"96", X"96", X"96"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"91", X"91", X"91"), (X"ED", X"ED", X"ED"), (X"92", X"92", X"92"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"96", X"96", X"96"), (X"EB", X"EB", X"EB"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"9A", X"9A", X"9A"), (X"E6", X"E6", X"E6"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"9F", X"9F", X"9F"), (X"E2", X"E2", X"E2"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"A3", X"A3", X"A3"), (X"DD", X"DD", X"DD"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"A9", X"A9", X"A9"), (X"D7", X"D7", X"D7"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"B0", X"B0", X"B0"), (X"D1", X"D1", X"D1"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"B6", X"B6", X"B6"), (X"CA", X"CA", X"CA"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"90", X"90", X"90"), (X"BD", X"BD", X"BD"), (X"8D", X"8D", X"8D"), (X"2B", X"2B", X"2B"), (X"2B", X"2B", X"2B"), (X"2B", X"2B", X"2B"), (X"2B", X"2B", X"2B"), (X"2B", X"2B", X"2B"), (X"2B", X"2B", X"2B"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"A7", X"A7", X"A7"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"A6", X"A6", X"A6"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"94", X"94", X"94"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"B9", X"B9", X"B9"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"80", X"80", X"80"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"CD", X"CD", X"CD"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FC", X"FC", X"FC"), (X"70", X"70", X"70"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"E0", X"E0", X"E0"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F5", X"F5", X"F5"), (X"63", X"63", X"63"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5C", X"5C", X"5C"), (X"F2", X"F2", X"F2"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"EB", X"EB", X"EB"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"69", X"69", X"69"), (X"F8", X"F8", X"F8"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"D7", X"D7", X"D7"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"76", X"76", X"76"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"C4", X"C4", X"C4"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"89", X"89", X"89"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"B0", X"B0", X"B0"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"5A", X"5A", X"5A"), (X"9D", X"9D", X"9D"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"75", X"75", X"75"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"59", X"59", X"59"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"93", X"93", X"93"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"3B", X"3B", X"3B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"B2", X"B2", X"B2"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FA", X"FA", X"FA"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"D0", X"D0", X"D0"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F0", X"F0", X"F0"), (X"0E", X"0E", X"0E"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"EA", X"EA", X"EA"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"E0", X"E0", X"E0"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"17", X"17", X"17"), (X"F5", X"F5", X"F5"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"C1", X"C1", X"C1"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2B", X"2B", X"2B"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"A3", X"A3", X"A3"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"85", X"85", X"85"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"75", X"75", X"75"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"59", X"59", X"59"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"93", X"93", X"93"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"3B", X"3B", X"3B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"B2", X"B2", X"B2"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FA", X"FA", X"FA"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"D0", X"D0", X"D0"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F0", X"F0", X"F0"), (X"0E", X"0E", X"0E"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"EA", X"EA", X"EA"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"E0", X"E0", X"E0"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"17", X"17", X"17"), (X"F5", X"F5", X"F5"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"C1", X"C1", X"C1"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2B", X"2B", X"2B"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"A3", X"A3", X"A3"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"85", X"85", X"85"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), 
	(X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"77", X"77", X"77"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"75", X"75", X"75"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"59", X"59", X"59"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"93", X"93", X"93"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"3B", X"3B", X"3B"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"B2", X"B2", X"B2"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FA", X"FA", X"FA"), (X"22", X"22", X"22"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"D0", X"D0", X"D0"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"F0", X"F0", X"F0"), (X"0E", X"0E", X"0E"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"03", X"03", X"03"), (X"EA", X"EA", X"EA"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"E0", X"E0", X"E0"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"17", X"17", X"17"), (X"F5", X"F5", X"F5"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"C1", X"C1", X"C1"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"2B", X"2B", X"2B"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"A3", X"A3", X"A3"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"49", X"49", X"49"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"85", X"85", X"85"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"00", X"00", X"00"), (X"67", X"67", X"67"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF"), (X"FF", X"FF", X"FF")
);

begin

	process(clk)
	begin
	if(rising_edge(clk)) then
		q <= rom(addr);
	end if;
	end process;

end rtl;
