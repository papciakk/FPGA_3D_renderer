use work.common.all;

package renderer_mesh is
	constant vertices : vertex_attr_arr_t(0 to 161) := (
		va(150, -258, -16383, 127, 127, 0), va(-4284, -258, -15759, 92, 127, 4), va(-1217, 4066, -15759, 116, 159, 4), va(-8380, -258, -13938, 60, 127, 18), va(-5720, 4115, -14654, 80, 160, 13), va(-2486, 8060, -13938, 106, 190, 18), va(-11829, -258, -11052, 33, 127, 41), va(-9878, 4147, -12130, 48, 161, 33), va(-7033, 8158, -12130, 70, 191, 33), va(-3550, 11424, -11052, 97, 216, 41), va(-14367, -258, -7327, 13, 127, 70), 
		va(-13200, 4066, -8284, 22, 160, 62), va(-11017, 8060, -8615, 39, 190, 60), va(-7985, 11424, -8284, 63, 216, 62), va(-4335, 13896, -7327, 91, 235, 70), va(3738, 2412, -15759, 154, 147, 4), va(2394, 6818, -14654, 144, 181, 13), va(7053, 4885, -13938, 180, 166, 18), va(1139, 10878, -12130, 135, 212, 33), va(5740, 9347, -12130, 170, 200, 33), va(9844, 6962, -11052, 202, 182, 41), 
		va(37, 14096, -8284, 126, 236, 62), va(4417, 13204, -8615, 160, 229, 60), va(8472, 11284, -8284, 191, 215, 62), va(11897, 8490, -7327, 218, 193, 70), va(3738, -2930, -15759, 154, 106, 4), va(7408, -258, -14654, 184, 127, 13), va(7053, -5399, -13938, 180, 87, 18), va(10788, 2220, -12130, 210, 145, 33), va(10788, -2738, -12130, 210, 108, 33), va(9844, -7479, -11052, 202, 71, 41), 
		va(13432, 4287, -8284, 230, 161, 62), va(13957, -258, -8615, 235, 127, 60), va(13432, -4804, -8284, 230, 92, 62), va(11897, -9008, -7327, 218, 60, 70), va(-1217, -4584, -15759, 116, 94, 4), va(2394, -7336, -14654, 144, 72, 13), va(-2486, -8577, -13938, 106, 63, 18), va(5740, -9864, -12130, 170, 53, 33), va(1139, -11396, -12130, 135, 41, 33), va(-3550, -11941, -11052, 97, 37, 41), 
		va(8472, -11802, -8284, 191, 38, 62), va(4417, -13721, -8615, 160, 24, 60), va(37, -14613, -8284, 126, 17, 62), va(-4335, -14414, -7327, 91, 18, 70), va(-5720, -4633, -14654, 80, 93, 13), va(-7033, -8675, -12130, 70, 62, 33), va(-9878, -4661, -12130, 48, 92, 33), va(-7985, -11941, -8284, 63, 37, 62), va(-11017, -8577, -8615, 39, 63, 60), va(-13200, -4584, -8284, 22, 93, 62), 
		va(-15417, -2930, -3808, 5, 106, 97), va(-15417, 2412, -3808, 5, 147, 97), va(-15284, -5399, 0, 6, 87, 127), va(-16079, -258, 0, 0, 127, 127), va(-15284, 4885, 0, 6, 166, 127), va(-13978, -7479, 3808, 16, 72, 156), va(-15356, -2738, 4180, 5, 108, 159), va(-15356, 2220, 4180, 5, 145, 159), va(-13978, 6962, 3808, 16, 181, 156), va(-11593, -9008, 7327, 35, 60, 183), 
		va(-13128, -4804, 8284, 23, 92, 191), va(-13654, -258, 8615, 18, 127, 193), va(-13128, 4287, 8284, 23, 161, 191), va(-11593, 8490, 7327, 35, 193, 183), va(-7139, 14096, -3808, 69, 236, 97), va(-2179, 15746, -3808, 108, 249, 97), va(-9390, 13204, 0, 52, 229, 127), va(-4864, 15568, 0, 87, 247, 127), va(150, 16383, 0, 127, 254, 127), va(-10911, 11284, 3808, 40, 215, 156), 
		va(-6941, 14092, 4180, 71, 236, 159), va(-2339, 15627, 4180, 107, 248, 159), va(2483, 15746, 3808, 145, 249, 156), va(-8172, 11284, 8284, 62, 215, 191), va(-4113, 13204, 8615, 93, 229, 193), va(266, 14096, 8284, 127, 236, 191), va(4638, 13896, 7327, 162, 235, 183), va(11215, 11284, -3808, 213, 215, 97), va(14278, 6962, -3808, 237, 181, 97), va(9690, 13204, 0, 201, 229, 127), 
		va(13282, 9522, 0, 229, 201, 127), va(15588, 4885, 0, 247, 166, 127), va(7442, 14096, 3808, 184, 236, 156), va(11273, 11092, 4180, 214, 213, 159), va(14118, 7077, 4180, 236, 183, 159), va(15721, 2412, 3808, 248, 147, 156), va(8288, 11424, 8284, 190, 216, 191), va(11321, 8060, 8615, 214, 190, 193), va(13504, 4066, 8284, 231, 160, 191), va(14667, -258, 7327, 240, 127, 183), 
		va(14278, -7479, -3808, 237, 72, 97), va(11215, -11802, -3808, 213, 38, 97), va(15588, -5399, 0, 247, 87, 127), va(13282, -10039, 0, 229, 52, 127), va(9690, -13721, 0, 201, 24, 127), va(15721, -2930, 3808, 248, 106, 156), va(14118, -7595, 4180, 236, 70, 159), va(11273, -11609, 4180, 214, 40, 159), va(7442, -14613, 3808, 184, 17, 156), va(13504, -4584, 8284, 231, 93, 191), 
		va(11321, -8577, 8615, 214, 63, 193), va(8288, -11941, 8284, 190, 37, 191), va(4638, -14414, 7327, 162, 18, 183), va(-2179, -16264, -3808, 108, 4, 97), va(-7139, -14613, -3808, 69, 17, 97), va(150, -16897, 0, 127, 0, 127), va(-4864, -16082, 0, 87, 6, 127), va(-9390, -13721, 0, 52, 24, 127), va(2483, -16264, 3808, 145, 4, 156), va(-2339, -16145, 4180, 107, 5, 159), 
		va(-6941, -14610, 4180, 71, 17, 159), va(-10911, -11802, 3808, 40, 38, 156), va(266, -14613, 8284, 127, 17, 191), va(-4113, -13721, 8615, 93, 24, 193), va(-8172, -11802, 8284, 62, 38, 191), va(-12978, 9522, 0, 24, 201, 126), va(-10973, 11092, -4180, 39, 213, 94), va(-13814, 7077, -4180, 17, 183, 94), va(5167, 15568, 0, 166, 247, 126), va(7244, 14092, -4180, 182, 236, 94), 
		va(2643, 15627, -4180, 146, 248, 94), va(16383, -258, 0, 253, 127, 126), va(15656, -2738, -4180, 248, 108, 94), va(15656, 2220, -4180, 248, 145, 94), va(5167, -16082, 0, 166, 6, 126), va(2643, -16145, -4180, 146, 5, 94), va(7244, -14610, -4180, 182, 17, 94), va(-12978, -10039, 0, 24, 52, 126), va(-13814, -7595, -4180, 17, 70, 94), va(-10973, -11609, -4180, 39, 40, 94), 
		va(150, -258, 16383, 127, 127, 254), va(1521, 4066, 15759, 137, 159, 249), va(-3438, 2412, 15759, 99, 147, 249), va(2786, 8060, 13938, 147, 190, 235), va(-2090, 6818, 14654, 109, 181, 240), va(-6753, 4885, 13938, 73, 166, 235), va(3854, 11424, 11052, 156, 216, 212), va(-835, 10878, 12130, 118, 212, 220), va(-5437, 9347, 12130, 83, 200, 220), va(-9540, 6962, 11052, 51, 182, 212), 
		va(4587, -258, 15759, 161, 127, 249), va(8684, -258, 13938, 193, 127, 235), va(6023, 4115, 14654, 173, 160, 240), va(12132, -258, 11052, 220, 127, 212), va(10178, 4147, 12130, 205, 161, 220), va(7337, 8158, 12130, 183, 191, 220), va(1521, -4584, 15759, 137, 94, 249), va(2786, -8577, 13938, 147, 63, 235), va(6023, -4633, 14654, 173, 93, 240), va(3854, -11941, 11052, 156, 37, 212), 
		va(7337, -8675, 12130, 183, 62, 220), va(10178, -4661, 12130, 205, 92, 220), va(-3438, -2930, 15759, 99, 106, 249), va(-6753, -5399, 13938, 73, 87, 235), va(-2090, -7336, 14654, 109, 72, 240), va(-9540, -7479, 11052, 51, 71, 212), va(-5437, -9864, 12130, 83, 53, 220), va(-835, -11396, 12130, 118, 41, 220), va(-7108, -258, 14654, 69, 127, 240), va(-10488, 2220, 12130, 43, 145, 220), 
		va(-10488, -2738, 12130, 43, 108, 220)
	);

	constant indices : indices_arr_t(0 to 319) := (
		idx(0, 1, 2), idx(1, 3, 4), 
		idx(1, 4, 2), idx(2, 4, 5), idx(3, 6, 7), idx(3, 7, 4), idx(4, 7, 8), idx(4, 8, 5), idx(5, 8, 9), idx(6, 10, 11), idx(6, 11, 7), idx(7, 11, 12), 
		idx(7, 12, 8), idx(8, 12, 13), idx(8, 13, 9), idx(9, 13, 14), idx(0, 2, 15), idx(2, 5, 16), idx(2, 16, 15), idx(15, 16, 17), idx(5, 9, 18), idx(5, 18, 16), 
		idx(16, 18, 19), idx(16, 19, 17), idx(17, 19, 20), idx(9, 14, 21), idx(9, 21, 18), idx(18, 21, 22), idx(18, 22, 19), idx(19, 22, 23), idx(19, 23, 20), idx(20, 23, 24), 
		idx(0, 15, 25), idx(15, 17, 26), idx(15, 26, 25), idx(25, 26, 27), idx(17, 20, 28), idx(17, 28, 26), idx(26, 28, 29), idx(26, 29, 27), idx(27, 29, 30), idx(20, 24, 31), 
		idx(20, 31, 28), idx(28, 31, 32), idx(28, 32, 29), idx(29, 32, 33), idx(29, 33, 30), idx(30, 33, 34), idx(0, 25, 35), idx(25, 27, 36), idx(25, 36, 35), idx(35, 36, 37), 
		idx(27, 30, 38), idx(27, 38, 36), idx(36, 38, 39), idx(36, 39, 37), idx(37, 39, 40), idx(30, 34, 41), idx(30, 41, 38), idx(38, 41, 42), idx(38, 42, 39), idx(39, 42, 43), 
		idx(39, 43, 40), idx(40, 43, 44), idx(0, 35, 1), idx(35, 37, 45), idx(35, 45, 1), idx(1, 45, 3), idx(37, 40, 46), idx(37, 46, 45), idx(45, 46, 47), idx(45, 47, 3), 
		idx(3, 47, 6), idx(40, 44, 48), idx(40, 48, 46), idx(46, 48, 49), idx(46, 49, 47), idx(47, 49, 50), idx(47, 50, 6), idx(6, 50, 10), idx(10, 51, 52), idx(51, 53, 54), 
		idx(51, 54, 52), idx(52, 54, 55), idx(53, 56, 57), idx(53, 57, 54), idx(54, 57, 58), idx(54, 58, 55), idx(55, 58, 59), idx(56, 60, 61), idx(56, 61, 57), idx(57, 61, 62), 
		idx(57, 62, 58), idx(58, 62, 63), idx(58, 63, 59), idx(59, 63, 64), idx(14, 65, 66), idx(65, 67, 68), idx(65, 68, 66), idx(66, 68, 69), idx(67, 70, 71), idx(67, 71, 68), 
		idx(68, 71, 72), idx(68, 72, 69), idx(69, 72, 73), idx(70, 64, 74), idx(70, 74, 71), idx(71, 74, 75), idx(71, 75, 72), idx(72, 75, 76), idx(72, 76, 73), idx(73, 76, 77), 
		idx(24, 78, 79), idx(78, 80, 81), idx(78, 81, 79), idx(79, 81, 82), idx(80, 83, 84), idx(80, 84, 81), idx(81, 84, 85), idx(81, 85, 82), idx(82, 85, 86), idx(83, 77, 87), 
		idx(83, 87, 84), idx(84, 87, 88), idx(84, 88, 85), idx(85, 88, 89), idx(85, 89, 86), idx(86, 89, 90), idx(34, 91, 92), idx(91, 93, 94), idx(91, 94, 92), idx(92, 94, 95), 
		idx(93, 96, 97), idx(93, 97, 94), idx(94, 97, 98), idx(94, 98, 95), idx(95, 98, 99), idx(96, 90, 100), idx(96, 100, 97), idx(97, 100, 101), idx(97, 101, 98), idx(98, 101, 102), 
		idx(98, 102, 99), idx(99, 102, 103), idx(44, 104, 105), idx(104, 106, 107), idx(104, 107, 105), idx(105, 107, 108), idx(106, 109, 110), idx(106, 110, 107), idx(107, 110, 111), idx(107, 111, 108), 
		idx(108, 111, 112), idx(109, 103, 113), idx(109, 113, 110), idx(110, 113, 114), idx(110, 114, 111), idx(111, 114, 115), idx(111, 115, 112), idx(112, 115, 60), idx(64, 70, 59), idx(70, 67, 116), 
		idx(70, 116, 59), idx(59, 116, 55), idx(67, 65, 117), idx(67, 117, 116), idx(116, 117, 118), idx(116, 118, 55), idx(55, 118, 52), idx(65, 14, 13), idx(65, 13, 117), idx(117, 13, 12), 
		idx(117, 12, 118), idx(118, 12, 11), idx(118, 11, 52), idx(52, 11, 10), idx(77, 83, 73), idx(83, 80, 119), idx(83, 119, 73), idx(73, 119, 69), idx(80, 78, 120), idx(80, 120, 119), 
		idx(119, 120, 121), idx(119, 121, 69), idx(69, 121, 66), idx(78, 24, 23), idx(78, 23, 120), idx(120, 23, 22), idx(120, 22, 121), idx(121, 22, 21), idx(121, 21, 66), idx(66, 21, 14), 
		idx(90, 96, 86), idx(96, 93, 122), idx(96, 122, 86), idx(86, 122, 82), idx(93, 91, 123), idx(93, 123, 122), idx(122, 123, 124), idx(122, 124, 82), idx(82, 124, 79), idx(91, 34, 33), 
		idx(91, 33, 123), idx(123, 33, 32), idx(123, 32, 124), idx(124, 32, 31), idx(124, 31, 79), idx(79, 31, 24), idx(103, 109, 99), idx(109, 106, 125), idx(109, 125, 99), idx(99, 125, 95), 
		idx(106, 104, 126), idx(106, 126, 125), idx(125, 126, 127), idx(125, 127, 95), idx(95, 127, 92), idx(104, 44, 43), idx(104, 43, 126), idx(126, 43, 42), idx(126, 42, 127), idx(127, 42, 41), 
		idx(127, 41, 92), idx(92, 41, 34), idx(60, 56, 112), idx(56, 53, 128), idx(56, 128, 112), idx(112, 128, 108), idx(53, 51, 129), idx(53, 129, 128), idx(128, 129, 130), idx(128, 130, 108), 
		idx(108, 130, 105), idx(51, 10, 50), idx(51, 50, 129), idx(129, 50, 49), idx(129, 49, 130), idx(130, 49, 48), idx(130, 48, 105), idx(105, 48, 44), idx(131, 132, 133), idx(132, 134, 135), 
		idx(132, 135, 133), idx(133, 135, 136), idx(134, 137, 138), idx(134, 138, 135), idx(135, 138, 139), idx(135, 139, 136), idx(136, 139, 140), idx(137, 77, 76), idx(137, 76, 138), idx(138, 76, 75), 
		idx(138, 75, 139), idx(139, 75, 74), idx(139, 74, 140), idx(140, 74, 64), idx(131, 141, 132), idx(141, 142, 143), idx(141, 143, 132), idx(132, 143, 134), idx(142, 144, 145), idx(142, 145, 143), 
		idx(143, 145, 146), idx(143, 146, 134), idx(134, 146, 137), idx(144, 90, 89), idx(144, 89, 145), idx(145, 89, 88), idx(145, 88, 146), idx(146, 88, 87), idx(146, 87, 137), idx(137, 87, 77), 
		idx(131, 147, 141), idx(147, 148, 149), idx(147, 149, 141), idx(141, 149, 142), idx(148, 150, 151), idx(148, 151, 149), idx(149, 151, 152), idx(149, 152, 142), idx(142, 152, 144), idx(150, 103, 102), 
		idx(150, 102, 151), idx(151, 102, 101), idx(151, 101, 152), idx(152, 101, 100), idx(152, 100, 144), idx(144, 100, 90), idx(131, 153, 147), idx(153, 154, 155), idx(153, 155, 147), idx(147, 155, 148), 
		idx(154, 156, 157), idx(154, 157, 155), idx(155, 157, 158), idx(155, 158, 148), idx(148, 158, 150), idx(156, 60, 115), idx(156, 115, 157), idx(157, 115, 114), idx(157, 114, 158), idx(158, 114, 113), 
		idx(158, 113, 150), idx(150, 113, 103), idx(131, 133, 153), idx(133, 136, 159), idx(133, 159, 153), idx(153, 159, 154), idx(136, 140, 160), idx(136, 160, 159), idx(159, 160, 161), idx(159, 161, 154), 
		idx(154, 161, 156), idx(140, 64, 63), idx(140, 63, 160), idx(160, 63, 62), idx(160, 62, 161), idx(161, 62, 61), idx(161, 61, 156), idx(156, 61, 60)
	);

end package renderer_mesh;
