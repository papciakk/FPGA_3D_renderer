use work.definitions.all;

package mesh is
	constant vertices : vertex_attr_arr_t(0 to 45) := (
		va(0, 0, 29929, 0, 0, 32767), va(0, 16181, 25178, 0, 18835, 26813), va(-8748, 13612, 25178, -10183, 15845, 26813), 
		va(-14718, 6721, 25178, -17133, 7824, 26813), va(-16016, -2302, 25178, -18643, -2681, 26813), va(-12228, -10596, 25178, -14235, -12334, 26813), 
		va(-4558, -15525, 25178, -5306, -18072, 26813), va(4558, -15525, 25178, 5306, -18072, 26813), va(12228, -10596, 25178, 14235, -12334, 26813), 
		va(16016, -2302, 25178, 18643, -2681, 26813), va(14718, 6721, 25178, 17133, 7824, 26813), va(8748, 13612, 25178, 10183, 15845, 26813), 
		va(0, 27224, 12433, 0, 30068, 13022), va(-14718, 22903, 12433, -16256, 25295, 13022), va(-24764, 11309, 12433, -27351, 12491, 13022), 
		va(-26947, -3874, 12433, -29762, -4279, 13022), va(-20575, -17828, 12433, -22724, -19691, 13022), va(-7670, -26122, 12433, -8471, -28850, 13022), 
		va(7670, -26122, 12433, 8471, -28850, 13022), va(20575, -17828, 12433, 22724, -19691, 13022), va(26947, -3874, 12433, 29762, -4279, 13022), 
		va(24764, 11309, 12433, 27351, 12491, 13022), va(14718, 22903, 12433, 16256, 25295, 13022), va(0, 29625, -4259, 0, 32464, -4446), 
		va(-16016, 24922, -4259, -17551, 27310, -4446), va(-26947, 12306, -4259, -29530, 13486, -4446), va(-29323, -4216, -4259, -32134, -4620, -4446), 
		va(-22389, -19400, -4259, -24535, -21259, -4446), va(-8346, -28425, -4259, -9146, -31149, -4446), va(8346, -28425, -4259, 9146, -31149, -4446), 
		va(22389, -19400, -4259, 24535, -21259, -4446), va(29323, -4216, -4259, 32134, -4620, -4446), va(26947, 12306, -4259, 29530, 13486, -4446), 
		va(16016, 24922, -4259, 17551, 27310, -4446), va(0, 22619, -19599, 0, 24118, -22181), va(-12228, 19028, -19599, -13039, 20289, -22181), 
		va(-20575, 9396, -19599, -21938, 10019, -22181), va(-22389, -3219, -19599, -23872, -3432, -22181), va(-17094, -14812, -19599, -18227, -15794, -22181), 
		va(-6372, -21703, -19599, -6795, -23141, -22181), va(6372, -21703, -19599, 6795, -23141, -22181), va(17094, -14812, -19599, 18227, -15794, -22181), 
		va(22389, -3219, -19599, 23872, -3432, -22181), va(20575, 9396, -19599, 21938, 10019, -22181), va(12228, 19028, -19599, 13039, 20289, -22181), 
		va(0, 0, -29929, 0, 0, -32767)
	);

	constant indices : indices_arr_t(0 to 87) := (
		idx(0, 1, 2), idx(0, 2, 3), idx(0, 3, 4), idx(0, 4, 5), idx(0, 5, 6), 
		idx(0, 6, 7), idx(0, 7, 8), idx(0, 8, 9), idx(0, 9, 10), idx(0, 10, 11), 
		idx(0, 11, 1), idx(1, 12, 13), idx(1, 13, 2), idx(2, 13, 14), idx(2, 14, 3), 
		idx(3, 14, 15), idx(3, 15, 4), idx(4, 15, 16), idx(4, 16, 5), idx(5, 16, 17), 
		idx(5, 17, 6), idx(6, 17, 18), idx(6, 18, 7), idx(7, 18, 19), idx(7, 19, 8), 
		idx(8, 19, 20), idx(8, 20, 9), idx(9, 20, 21), idx(9, 21, 10), idx(10, 21, 22), 
		idx(10, 22, 11), idx(11, 22, 12), idx(11, 12, 1), idx(12, 23, 24), idx(12, 24, 13), 
		idx(13, 24, 25), idx(13, 25, 14), idx(14, 25, 26), idx(14, 26, 15), idx(15, 26, 27), 
		idx(15, 27, 16), idx(16, 27, 28), idx(16, 28, 17), idx(17, 28, 29), idx(17, 29, 18), 
		idx(18, 29, 30), idx(18, 30, 19), idx(19, 30, 31), idx(19, 31, 20), idx(20, 31, 32), 
		idx(20, 32, 21), idx(21, 32, 33), idx(21, 33, 22), idx(22, 33, 23), idx(22, 23, 12), 
		idx(23, 34, 35), idx(23, 35, 24), idx(24, 35, 36), idx(24, 36, 25), idx(25, 36, 37), 
		idx(25, 37, 26), idx(26, 37, 38), idx(26, 38, 27), idx(27, 38, 39), idx(27, 39, 28), 
		idx(28, 39, 40), idx(28, 40, 29), idx(29, 40, 41), idx(29, 41, 30), idx(30, 41, 42), 
		idx(30, 42, 31), idx(31, 42, 43), idx(31, 43, 32), idx(32, 43, 44), idx(32, 44, 33), 
		idx(33, 44, 34), idx(33, 34, 23), idx(45, 35, 34), idx(45, 36, 35), idx(45, 37, 36), 
		idx(45, 38, 37), idx(45, 39, 38), idx(45, 40, 39), idx(45, 41, 40), idx(45, 42, 41), 
		idx(45, 43, 42), idx(45, 44, 43), idx(45, 34, 44)
	);

end package;
